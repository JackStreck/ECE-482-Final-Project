* ==========================================================
* C2MOS REGISTER — PARAMETRIC SIZING + FUNCTIONALITY TEST
* ==========================================================

.lib '/class/ece482/gpdk045_mos' TT

.TEMP 25
.OPTION POST

* ----------------------------------------------------------
* SIZING PARAMETERS (EDIT THESE TO TUNE THE REGISTER)
* ----------------------------------------------------------
* Base “unit” sizes
.param wn_unit = 120n
.param wp_unit = 240n

* Global scaling factor (you can also .step this)
.param k_size = 1.0

* Individual device groups (you can tweak ratios here)
.param wn_d   = k_size * wn_unit
.param wn_clk = k_size * wn_unit
.param wn_q   = k_size * wn_unit
.param wn_rst = k_size * wn_unit

.param wp_d   = k_size * wp_unit
.param wp_clk = k_size * wp_unit
.param wp_q   = k_size * wp_unit

* ----------------------------------------------------------
* SUPPLIES
* ----------------------------------------------------------
VDD   vdd   0  1.1
VSS   vss   0  0

* ----------------------------------------------------------
* INPUT STIMULI
* ----------------------------------------------------------
* Clock: 0–1.1 V, 4 ns period (2 ns high, 2 ns low)
VCLK      clk      0  PULSE(0 1.1 0 20p 20p 2n 4n)
* Complement clock (ideal, for C2MOS; duty matches)
VCLK_BAR  clk_bar  0  PULSE(1.1 0 0 20p 20p 2n 4n)

* Data input: changes slower than clock so you can see sampling
* Example: D low first 8 ns, then high 8–16 ns, then low again
VD        d        0  PWL(0n 0   7.9n 0   8n 1.1   15.9n 1.1   16n 0   40n 0)

* Asynchronous reset (assume active-high, clears Q=0 initially)
* High from 0–3 ns, then low (released)
VRST      rst      0  PWL(0n 1.1   3n 1.1   3.1n 0   40n 0)

* ----------------------------------------------------------
* EXTRACTED C2MOS REGISTER DEVICES
* (Your giant layout-extracted blob, unchanged except for params)
* ----------------------------------------------------------

** Library name: test2
** Cell name: C2MOS_register
** View name: schematic

mpm3 net17 x vdd vdd g45p1svt L=45e-9 W=wp_q AD='wp_q/ceil((wp_q-5e-12)/10e-6)<119.5e-9?(floor(ceil((wp_q-5e-12)/10e-6)/2.0)*(14.4e-15+(wp_q/ceil((wp_q-5e-12)/10e-6))*100e-9)+(ceil((wp_q-5e-12)/10e-6)/2-floor(ceil((wp_q-5e-12)/10e-6)/2)!=0?14.4e-15+(wp_q/ceil((wp_q-5e-12)/10e-6))*50e-9:0))/1:(floor(ceil((wp_q-5e-12)/10e-6)/2.0)*(110e-9*(wp_q/ceil((wp_q-5e-12)/10e-6)))+(ceil((wp_q-5e-12)/10e-6)/2-floor(ceil((wp_q-5e-12)/10e-6)/2)!=0?140e-9*(wp_q/ceil((wp_q-5e-12)/10e-6)):0))/1' AS='wp_q/ceil((wp_q-5e-12)/10e-6)<119.5e-9?(((14.4e-15+(wp_q/ceil((wp_q-5e-12)/10e-6))*50e-9)+floor((ceil((wp_q-5e-12)/10e-6)-1)/2.0)*(14.4e-15+(wp_q/ceil((wp_q-5e-12)/10e-6))*100e-9))+(ceil((wp_q-5e-12)/10e-6)/2-floor(ceil((wp_q-5e-12)/10e-6)/2)==0?14.4e-15+(wp_q/ceil((wp_q-5e-12)/10e-6))*50e-9:0))/1:((140e-9*(wp_q/ceil((wp_q-5e-12)/10e-6))+floor((ceil((wp_q-5e-12)/10e-6)-1)/2.0)*(110e-9*(wp_q/ceil((wp_q-5e-12)/10e-6))))+(ceil((wp_q-5e-12)/10e-6)/2-floor(ceil((wp_q-5e-12)/10e-6)/2)==0?140e-9*(wp_q/ceil((wp_q-5e-12)/10e-6)):0))/1'
+PD='wp_q/ceil((wp_q-5e-12)/10e-6)<119.5e-9?(floor(ceil((wp_q-5e-12)/10e-6)/2.0)*680e-9+(ceil((wp_q-5e-12)/10e-6)/2-floor(ceil((wp_q-5e-12)/10e-6)/2)!=0?580e-9:0))/1:(floor(ceil((wp_q-5e-12)/10e-6)/2.0)*(220e-9+2*(wp_q/ceil((wp_q-5e-12)/10e-6)))+(ceil((wp_q-5e-12)/10e-6)/2-floor(ceil((wp_q-5e-12)/10e-6)/2)!=0?280e-9+2*(wp_q/ceil((wp_q-5e-12)/10e-6)):0))/1' PS='wp_q/ceil((wp_q-5e-12)/10e-6)<119.5e-9?((580e-9+floor((ceil((wp_q-5e-12)/10e-6)-1)/2.0)*680e-9)+(ceil((wp_q-5e-12)/10e-6)/2-floor(ceil((wp_q-5e-12)/10e-6)/2)==0?580e-9:0))/1:(((280e-9+2*(wp_q/ceil((wp_q-5e-12)/10e-6)))+floor((ceil((wp_q-5e-12)/10e-6)-1)/2.0)*(220e-9+2*(wp_q/ceil((wp_q-5e-12)/10e-6))))+(ceil((wp_q-5e-12)/10e-6)/2-floor(ceil((wp_q-5e-12)/10e-6)/2)==0?280e-9+2*(wp_q/ceil((wp_q-5e-12)/10e-6)):0))/1'
+NRD='wp_q/ceil((wp_q-5e-12)/10e-6)<119.5e-9?(floor(ceil((wp_q-5e-12)/10e-6)/2.0)*(14.4e-15+(wp_q/ceil((wp_q-5e-12)/10e-6))*100e-9)+(ceil((wp_q-5e-12)/10e-6)/2-floor(ceil((wp_q-5e-12)/10e-6)/2)!=0?14.4e-15+(wp_q/ceil((wp_q-5e-12)/10e-6))*50e-9:0))/1:((floor(ceil((wp_q-5e-12)/10e-6)/2.0)*(110e-9*(wp_q/ceil((wp_q-5e-12)/10e-6)))+(ceil((wp_q-5e-12)/10e-6)/2-floor(ceil((wp_q-5e-12)/10e-6)/2)!=0?140e-9*(wp_q/ceil((wp_q-5e-12)/10e-6)):0))/1)/((((wp_q/ceil((wp_q-5e-12)/10e-6))*ceil((wp_q-5e-12)/10e-6))*(wp_q/ceil((wp_q-5e-12)/10e-6)))*ceil((wp_q-5e-12)/10e-6))'
+NRS='wp_q/ceil((wp_q-5e-12)/10e-6)<119.5e-9?(((14.4e-15+(wp_q/ceil((wp_q-5e-12)/10e-6))*50e-9)+floor((ceil((wp_q-5e-12)/10e-6)-1)/2.0)*(14.4e-15+(wp_q/ceil((wp_q-5e-12)/10e-6))*100e-9))+(ceil((wp_q-5e-12)/10e-6)/2-floor(ceil((wp_q-5e-12)/10e-6)/2)==0?14.4e-15+(wp_q/ceil((wp_q-5e-12)/10e-6))*50e-9:0))/1:(((140e-9*(wp_q/ceil((wp_q-5e-12)/10e-6))+floor((ceil((wp_q-5e-12)/10e-6)-1)/2.0)*(110e-9*(wp_q/ceil((wp_q-5e-12)/10e-6))))+(ceil((wp_q-5e-12)/10e-6)/2-floor(ceil((wp_q-5e-12)/10e-6)/2)==0?140e-9*(wp_q/ceil((wp_q-5e-12)/10e-6)):0))/1)/((((wp_q/ceil((wp_q-5e-12)/10e-6))*ceil((wp_q-5e-12)/10e-6))*(wp_q/ceil((wp_q-5e-12)/10e-6)))*ceil((wp_q-5e-12)/10e-6))' M=1

mpm2 q clk_bar net17 vdd g45p1svt L=45e-9 W=wp_clk AD='wp_clk/ceil((wp_clk-5e-12)/10e-6)<119.5e-9?(floor(ceil((wp_clk-5e-12)/10e-6)/2.0)*(14.4e-15+(wp_clk/ceil((wp_clk-5e-12)/10e-6))*100e-9)+(ceil((wp_clk-5e-12)/10e-6)/2-floor(ceil((wp_clk-5e-12)/10e-6)/2)!=0?14.4e-15+(wp_clk/ceil((wp_clk-5e-12)/10e-6))*50e-9:0))/1:(floor(ceil((wp_clk-5e-12)/10e-6)/2.0)*(110e-9*(wp_clk/ceil((wp_clk-5e-12)/10e-6)))+(ceil((wp_clk-5e-12)/10e-6)/2-floor(ceil((wp_clk-5e-12)/10e-6)/2)!=0?140e-9*(wp_clk/ceil((wp_clk-5e-12)/10e-6)):0))/1'
+AS='wp_clk/ceil((wp_clk-5e-12)/10e-6)<119.5e-9?(((14.4e-15+(wp_clk/ceil((wp_clk-5e-12)/10e-6))*50e-9)+floor((ceil((wp_clk-5e-12)/10e-6)-1)/2.0)*(14.4e-15+(wp_clk/ceil((wp_clk-5e-12)/10e-6))*100e-9))+(ceil((wp_clk-5e-12)/10e-6)/2-floor(ceil((wp_clk-5e-12)/10e-6)/2)==0?14.4e-15+(wp_clk/ceil((wp_clk-5e-12)/10e-6))*50e-9:0))/1:((140e-9*(wp_clk/ceil((wp_clk-5e-12)/10e-6))+floor((ceil((wp_clk-5e-12)/10e-6)-1)/2.0)*(110e-9*(wp_clk/ceil((wp_clk-5e-12)/10e-6))))+(ceil((wp_clk-5e-12)/10e-6)/2-floor(ceil((wp_clk-5e-12)/10e-6)/2)==0?140e-9*(wp_clk/ceil((wp_clk-5e-12)/10e-6)):0))/1' PD='wp_clk/ceil((wp_clk-5e-12)/10e-6)<119.5e-9?(floor(ceil((wp_clk-5e-12)/10e-6)/2.0)*680e-9+(ceil((wp_clk-5e-12)/10e-6)/2-floor(ceil((wp_clk-5e-12)/10e-6)/2)!=0?580e-9:0))/1:(floor(ceil((wp_clk-5e-12)/10e-6)/2.0)*(220e-9+2*(wp_clk/ceil((wp_clk-5e-12)/10e-6)))+(ceil((wp_clk-5e-12)/10e-6)/2-floor(ceil((wp_clk-5e-12)/10e-6)/2)!=0?280e-9+2*(wp_clk/ceil((wp_clk-5e-12)/10e-6)):0))/1'
+PS='wp_clk/ceil((wp_clk-5e-12)/10e-6)<119.5e-9?((580e-9+floor((ceil((wp_clk-5e-12)/10e-6)-1)/2.0)*680e-9)+(ceil((wp_clk-5e-12)/10e-6)/2-floor(ceil((wp_clk-5e-12)/10e-6)/2)==0?580e-9:0))/1:(((280e-9+2*(wp_clk/ceil((wp_clk-5e-12)/10e-6)))+floor((ceil((wp_clk-5e-12)/10e-6)-1)/2.0)*(220e-9+2*(wp_clk/ceil((wp_clk-5e-12)/10e-6))))+(ceil((wp_clk-5e-12)/10e-6)/2-floor(ceil((wp_clk-5e-12)/10e-6)/2)==0?280e-9+2*(wp_clk/ceil((wp_clk-5e-12)/10e-6)):0))/1'
+NRD='wp_clk/ceil((wp_clk-5e-12)/10e-6)<119.5e-9?(floor(ceil((wp_clk-5e-12)/10e-6)/2.0)*(14.4e-15+(wp_clk/ceil((wp_clk-5e-12)/10e-6))*100e-9)+(ceil((wp_clk-5e-12)/10e-6)/2-floor(ceil((wp_clk-5e-12)/10e-6)/2)!=0?14.4e-15+(wp_clk/ceil((wp_clk-5e-12)/10e-6))*50e-9:0))/1:((floor(ceil((wp_clk-5e-12)/10e-6)/2.0)*(110e-9*(wp_clk/ceil((wp_clk-5e-12)/10e-6)))+(ceil((wp_clk-5e-12)/10e-6)/2-floor(ceil((wp_clk-5e-12)/10e-6)/2)!=0?140e-9*(wp_clk/ceil((wp_clk-5e-12)/10e-6)):0))/1)/((((wp_clk/ceil((wp_clk-5e-12)/10e-6))*ceil((wp_clk-5e-12)/10e-6))*(wp_clk/ceil((wp_clk-5e-12)/10e-6)))*ceil((wp_clk-5e-12)/10e-6))'
+NRS='wp_clk/ceil((wp_clk-5e-12)/10e-6)<119.5e-9?(((14.4e-15+(wp_clk/ceil((wp_clk-5e-12)/10e-6))*50e-9)+floor((ceil((wp_clk-5e-12)/10e-6)-1)/2.0)*(14.4e-15+(wp_clk/ceil((wp_clk-5e-12)/10e-6))*100e-9))+(ceil((wp_clk-5e-12)/10e-6)/2-floor(ceil((wp_clk-5e-12)/10e-6)/2)==0?14.4e-15+(wp_clk/ceil((wp_clk-5e-12)/10e-6))*50e-9:0))/1:(((140e-9*(wp_clk/ceil((wp_clk-5e-12)/10e-6))+floor((ceil((wp_clk-5e-12)/10e-6)-1)/2.0)*(110e-9*(wp_clk/ceil((wp_clk-5e-12)/10e-6))))+(ceil((wp_clk-5e-12)/10e-6)/2-floor(ceil((wp_clk-5e-12)/10e-6)/2)==0?140e-9*(wp_clk/ceil((wp_clk-5e-12)/10e-6)):0))/1)/((((wp_clk/ceil((wp_clk-5e-12)/10e-6))*ceil((wp_clk-5e-12)/10e-6))*(wp_clk/ceil((wp_clk-5e-12)/10e-6)))*ceil((wp_clk-5e-12)/10e-6))' M=1

mpm1 x clk net4 vdd g45p1svt L=45e-9 W=wp_clk AD='wp_clk/ceil((wp_clk-5e-12)/10e-6)<119.5e-9?(floor(ceil((wp_clk-5e-12)/10e-6)/2.0)*(14.4e-15+(wp_clk/ceil((wp_clk-5e-12)/10e-6))*100e-9)+(ceil((wp_clk-5e-12)/10e-6)/2-floor(ceil((wp_clk-5e-12)/10e-6)/2)!=0?14.4e-15+(wp_clk/ceil((wp_clk-5e-12)/10e-6))*50e-9:0))/1:(floor(ceil((wp_clk-5e-12)/10e-6)/2.0)*(110e-9*(wp_clk/ceil((wp_clk-5e-12)/10e-6)))+(ceil((wp_clk-5e-12)/10e-6)/2-floor(ceil((wp_clk-5e-12)/10e-6)/2)!=0?140e-9*(wp_clk/ceil((wp_clk-5e-12)/10e-6)):0))/1'
+AS='wp_clk/ceil((wp_clk-5e-12)/10e-6)<119.5e-9?(((14.4e-15+(wp_clk/ceil((wp_clk-5e-12)/10e-6))*50e-9)+floor((ceil((wp_clk-5e-12)/10e-6)-1)/2.0)*(14.4e-15+(wp_clk/ceil((wp_clk-5e-12)/10e-6))*100e-9))+(ceil((wp_clk-5e-12)/10e-6)/2-floor(ceil((wp_clk-5e-12)/10e-6)/2)==0?14.4e-15+(wp_clk/ceil((wp_clk-5e-12)/10e-6))*50e-9:0))/1:((140e-9*(wp_clk/ceil((wp_clk-5e-12)/10e-6))+floor((ceil((wp_clk-5e-12)/10e-6)-1)/2.0)*(110e-9*(wp_clk/ceil((wp_clk-5e-12)/10e-6))))+(ceil((wp_clk-5e-12)/10e-6)/2-floor(ceil((wp_clk-5e-12)/10e-6)/2)==0?140e-9*(wp_clk/ceil((wp_clk-5e-12)/10e-6)):0))/1' PD='wp_clk/ceil((wp_clk-5e-12)/10e-6)<119.5e-9?(floor(ceil((wp_clk-5e-12)/10e-6)/2.0)*680e-9+(ceil((wp_clk-5e-12)/10e-6)/2-floor(ceil((wp_clk-5e-12)/10e-6)/2)!=0?580e-9:0))/1:(floor(ceil((wp_clk-5e-12)/10e-6)/2.0)*(220e-9+2*(wp_clk/ceil((wp_clk-5e-12)/10e-6)))+(ceil((wp_clk-5e-12)/10e-6)/2-floor(ceil((wp_clk-5e-12)/10e-6)/2)!=0?280e-9+2*(wp_clk/ceil((wp_clk-5e-12)/10e-6)):0))/1'
+PS='wp_clk/ceil((wp_clk-5e-12)/10e-6)<119.5e-9?((580e-9+floor((ceil((wp_clk-5e-12)/10e-6)-1)/2.0)*680e-9)+(ceil((wp_clk-5e-12)/10e-6)/2-floor(ceil((wp_clk-5e-12)/10e-6)/2)==0?580e-9:0))/1:(((280e-9+2*(wp_clk/ceil((wp_clk-5e-12)/10e-6)))+floor((ceil((wp_clk-5e-12)/10e-6)-1)/2.0)*(220e-9+2*(wp_clk/ceil((wp_clk-5e-12)/10e-6))))+(ceil((wp_clk-5e-12)/10e-6)/2-floor(ceil((wp_clk-5e-12)/10e-6)/2)==0?280e-9+2*(wp_clk/ceil((wp_clk-5e-12)/10e-6)):0))/1'
+NRD='wp_clk/ceil((wp_clk-5e-12)/10e-6)<119.5e-9?(floor(ceil((wp_clk-5e-12)/10e-6)/2.0)*(14.4e-15+(wp_clk/ceil((wp_clk-5e-12)/10e-6))*100e-9)+(ceil((wp_clk-5e-12)/10e-6)/2-floor(ceil((wp_clk-5e-12)/10e-6)/2)!=0?14.4e-15+(wp_clk/ceil((wp_clk-5e-12)/10e-6))*50e-9:0))/1:((floor(ceil((wp_clk-5e-12)/10e-6)/2.0)*(110e-9*(wp_clk/ceil((wp_clk-5e-12)/10e-6)))+(ceil((wp_clk-5e-12)/10e-6)/2-floor(ceil((wp_clk-5e-12)/10e-6)/2)!=0?140e-9*(wp_clk/ceil((wp_clk-5e-12)/10e-6)):0))/1)/((((wp_clk/ceil((wp_clk-5e-12)/10e-6))*ceil((wp_clk-5e-12)/10e-6))*(wp_clk/ceil((wp_clk-5e-12)/10e-6)))*ceil((wp_clk-5e-12)/10e-6))'
+NRS='wp_clk/ceil((wp_clk-5e-12)/10e-6)<119.5e-9?(((14.4e-15+(wp_clk/ceil((wp_clk-5e-12)/10e-6))*50e-9)+floor((ceil((wp_clk-5e-12)/10e-6)-1)/2.0)*(14.4e-15+(wp_clk/ceil((wp_clk-5e-12)/10e-6))*100e-9))+(ceil((wp_clk-5e-12)/10e-6)/2-floor(ceil((wp_clk-5e-12)/10e-6)/2)==0?14.4e-15+(wp_clk/ceil((wp_clk-5e-12)/10e-6))*50e-9:0))/1:(((140e-9*(wp_clk/ceil((wp_clk-5e-12)/10e-6))+floor((ceil((wp_clk-5e-12)/10e-6)-1)/2.0)*(110e-9*(wp_clk/ceil((wp_clk-5e-12)/10e-6))))+(ceil((wp_clk-5e-12)/10e-6)/2-floor(ceil((wp_clk-5e-12)/10e-6)/2)==0?140e-9*(wp_clk/ceil((wp_clk-5e-12)/10e-6)):0))/1)/((((wp_clk/ceil((wp_clk-5e-12)/10e-6))*ceil((wp_clk-5e-12)/10e-6))*(wp_clk/ceil((wp_clk-5e-12)/10e-6)))*ceil((wp_clk-5e-12)/10e-6))' M=1

mpm0 net4 d vdd vdd g45p1svt L=45e-9 W=wp_d AD='wp_d/ceil((wp_d-5e-12)/10e-6)<119.5e-9?(floor(ceil((wp_d-5e-12)/10e-6)/2.0)*(14.4e-15+(wp_d/ceil((wp_d-5e-12)/10e-6))*100e-9)+(ceil((wp_d-5e-12)/10e-6)/2-floor(ceil((wp_d-5e-12)/10e-6)/2)!=0?14.4e-15+(wp_d/ceil((wp_d-5e-12)/10e-6))*50e-9:0))/1:(floor(ceil((wp_d-5e-12)/10e-6)/2.0)*(110e-9*(wp_d/ceil((wp_d-5e-12)/10e-6)))+(ceil((wp_d-5e-12)/10e-6)/2-floor(ceil((wp_d-5e-12)/10e-6)/2)!=0?140e-9*(wp_d/ceil((wp_d-5e-12)/10e-6)):0))/1' AS='wp_d/ceil((wp_d-5e-12)/10e-6)<119.5e-9?(((14.4e-15+(wp_d/ceil((wp_d-5e-12)/10e-6))*50e-9)+floor((ceil((wp_d-5e-12)/10e-6)-1)/2.0)*(14.4e-15+(wp_d/ceil((wp_d-5e-12)/10e-6))*100e-9))+(ceil((wp_d-5e-12)/10e-6)/2-floor(ceil((wp_d-5e-12)/10e-6)/2)==0?14.4e-15+(wp_d/ceil((wp_d-5e-12)/10e-6))*50e-9:0))/1:((140e-9*(wp_d/ceil((wp_d-5e-12)/10e-6))+floor((ceil((wp_d-5e-12)/10e-6)-1)/2.0)*(110e-9*(wp_d/ceil((wp_d-5e-12)/10e-6))))+(ceil((wp_d-5e-12)/10e-6)/2-floor(ceil((wp_d-5e-12)/10e-6)/2)==0?140e-9*(wp_d/ceil((wp_d-5e-12)/10e-6)):0))/1'
+PD='wp_d/ceil((wp_d-5e-12)/10e-6)<119.5e-9?(floor(ceil((wp_d-5e-12)/10e-6)/2.0)*680e-9+(ceil((wp_d-5e-12)/10e-6)/2-floor(ceil((wp_d-5e-12)/10e-6)/2)!=0?580e-9:0))/1:(floor(ceil((wp_d-5e-12)/10e-6)/2.0)*(220e-9+2*(wp_d/ceil((wp_d-5e-12)/10e-6)))+(ceil((wp_d-5e-12)/10e-6)/2-floor(ceil((wp_d-5e-12)/10e-6)/2)!=0?280e-9+2*(wp_d/ceil((wp_d-5e-12)/10e-6)):0))/1' PS='wp_d/ceil((wp_d-5e-12)/10e-6)<119.5e-9?((580e-9+floor((ceil((wp_d-5e-12)/10e-6)-1)/2.0)*680e-9)+(ceil((wp_d-5e-12)/10e-6)/2-floor(ceil((wp_d-5e-12)/10e-6)/2)==0?580e-9:0))/1:(((280e-9+2*(wp_d/ceil((wp_d-5e-12)/10e-6)))+floor((ceil((wp_d-5e-12)/10e-6)-1)/2.0)*(220e-9+2*(wp_d/ceil((wp_d-5e-12)/10e-6))))+(ceil((wp_d-5e-12)/10e-6)/2-floor(ceil((wp_d-5e-12)/10e-6)/2)==0?280e-9+2*(wp_d/ceil((wp_d-5e-12)/10e-6)):0))/1'
+NRD='wp_d/ceil((wp_d-5e-12)/10e-6)<119.5e-9?(floor(ceil((wp_d-5e-12)/10e-6)/2.0)*(14.4e-15+(wp_d/ceil((wp_d-5e-12)/10e-6))*100e-9)+(ceil((wp_d-5e-12)/10e-6)/2-floor(ceil((wp_d-5e-12)/10e-6)/2)!=0?14.4e-15+(wp_d/ceil((wp_d-5e-12)/10e-6))*50e-9:0))/1:((floor(ceil((wp_d-5e-12)/10e-6)/2.0)*(110e-9*(wp_d/ceil((wp_d-5e-12)/10e-6)))+(ceil((wp_d-5e-12)/10e-6)/2-floor(ceil((wp_d-5e-12)/10e-6)/2)!=0?140e-9*(wp_d/ceil((wp_d-5e-12)/10e-6)):0))/1)/((((wp_d/ceil((wp_d-5e-12)/10e-6))*ceil((wp_d-5e-12)/10e-6))*(wp_d/ceil((wp_d-5e-12)/10e-6)))*ceil((wp_d-5e-12)/10e-6))'
+NRS='wp_d/ceil((wp_d-5e-12)/10e-6)<119.5e-9?(((14.4e-15+(wp_d/ceil((wp_d-5e-12)/10e-6))*50e-9)+floor((ceil((wp_d-5e-12)/10e-6)-1)/2.0)*(14.4e-15+(wp_d/ceil((wp_d-5e-12)/10e-6))*100e-9))+(ceil((wp_d-5e-12)/10e-6)/2-floor(ceil((wp_d-5e-12)/10e-6)/2)==0?14.4e-15+(wp_d/ceil((wp_d-5e-12)/10e-6))*50e-9:0))/1:(((140e-9*(wp_d/ceil((wp_d-5e-12)/10e-6))+floor((ceil((wp_d-5e-12)/10e-6)-1)/2.0)*(110e-9*(wp_d/ceil((wp_d-5e-12)/10e-6))))+(ceil((wp_d-5e-12)/10e-6)/2-floor(ceil((wp_d-5e-12)/10e-6)/2)==0?140e-9*(wp_d/ceil((wp_d-5e-12)/10e-6)):0))/1)/((((wp_d/ceil((wp_d-5e-12)/10e-6))*ceil((wp_d-5e-12)/10e-6))*(wp_d/ceil((wp_d-5e-12)/10e-6)))*ceil((wp_d-5e-12)/10e-6))' M=1

mnm5 q rst vss vss g45n1svt L=45e-9 W=wn_rst AD='wn_rst/ceil((wn_rst-5e-12)/10e-6)<119.5e-9?(floor(ceil((wn_rst-5e-12)/10e-6)/2.0)*(14.4e-15+(wn_rst/ceil((wn_rst-5e-12)/10e-6))*100e-9)+(ceil((wn_rst-5e-12)/10e-6)/2-floor(ceil((wn_rst-5e-12)/10e-6)/2)!=0?14.4e-15+(wn_rst/ceil((wn_rst-5e-12)/10e-6))*50e-9:0))/1:(floor(ceil((wn_rst-5e-12)/10e-6)/2.0)*(110e-9*(wn_rst/ceil((wn_rst-5e-12)/10e-6)))+(ceil((wn_rst-5e-12)/10e-6)/2-floor(ceil((wn_rst-5e-12)/10e-6)/2)!=0?140e-9*(wn_rst/ceil((wn_rst-5e-12)/10e-6)):0))/1'
+AS='wn_rst/ceil((wn_rst-5e-12)/10e-6)<119.5e-9?(((14.4e-15+(wn_rst/ceil((wn_rst-5e-12)/10e-6))*50e-9)+floor((ceil((wn_rst-5e-12)/10e-6)-1)/2.0)*(14.4e-15+(wn_rst/ceil((wn_rst-5e-12)/10e-6))*100e-9))+(ceil((wn_rst-5e-12)/10e-6)/2-floor(ceil((wn_rst-5e-12)/10e-6)/2)==0?14.4e-15+(wn_rst/ceil((wn_rst-5e-12)/10e-6))*50e-9:0))/1:((140e-9*(wn_rst/ceil((wn_rst-5e-12)/10e-6))+floor((ceil((wn_rst-5e-12)/10e-6)-1)/2.0)*(110e-9*(wn_rst/ceil((wn_rst-5e-12)/10e-6))))+(ceil((wn_rst-5e-12)/10e-6)/2-floor(ceil((wn_rst-5e-12)/10e-6)/2)==0?140e-9*(wn_rst/ceil((wn_rst-5e-12)/10e-6)):0))/1' PD='wn_rst/ceil((wn_rst-5e-12)/10e-6)<119.5e-9?(floor(ceil((wn_rst-5e-12)/10e-6)/2.0)*680e-9+(ceil((wn_rst-5e-12)/10e-6)/2-floor(ceil((wn_rst-5e-12)/10e-6)/2)!=0?580e-9:0))/1:(floor(ceil((wn_rst-5e-12)/10e-6)/2.0)*(220e-9+2*(wn_rst/ceil((wn_rst-5e-12)/10e-6)))+(ceil((wn_rst-5e-12)/10e-6)/2-floor(ceil((wn_rst-5e-12)/10e-6)/2)!=0?280e-9+2*(wn_rst/ceil((wn_rst-5e-12)/10e-6)):0))/1'
+PS='wn_rst/ceil((wn_rst-5e-12)/10e-6)<119.5e-9?((580e-9+floor((ceil((wn_rst-5e-12)/10e-6)-1)/2.0)*680e-9)+(ceil((wn_rst-5e-12)/10e-6)/2-floor(ceil((wn_rst-5e-12)/10e-6)/2)==0?580e-9:0))/1:(((280e-9+2*(wn_rst/ceil((wn_rst-5e-12)/10e-6)))+floor((ceil((wn_rst-5e-12)/10e-6)-1)/2.0)*(220e-9+2*(wn_rst/ceil((wn_rst-5e-12)/10e-6))))+(ceil((wn_rst-5e-12)/10e-6)/2-floor(ceil((wn_rst-5e-12)/10e-6)/2)==0?280e-9+2*(wn_rst/ceil((wn_rst-5e-12)/10e-6)):0))/1'
+NRD='wn_rst/ceil((wn_rst-5e-12)/10e-6)<119.5e-9?(floor(ceil((wn_rst-5e-12)/10e-6)/2.0)*(14.4e-15+(wn_rst/ceil((wn_rst-5e-12)/10e-6))*100e-9)+(ceil((wn_rst-5e-12)/10e-6)/2-floor(ceil((wn_rst-5e-12)/10e-6)/2)!=0?14.4e-15+(wn_rst/ceil((wn_rst-5e-12)/10e-6))*50e-9:0))/1:((floor(ceil((wn_rst-5e-12)/10e-6)/2.0)*(110e-9*(wn_rst/ceil((wn_rst-5e-12)/10e-6)))+(ceil((wn_rst-5e-12)/10e-6)/2-floor(ceil((wn_rst-5e-12)/10e-6)/2)!=0?140e-9*(wn_rst/ceil((wn_rst-5e-12)/10e-6)):0))/1)/((((wn_rst/ceil((wn_rst-5e-12)/10e-6))*ceil((wn_rst-5e-12)/10e-6))*(wn_rst/ceil((wn_rst-5e-12)/10e-6)))*ceil((wn_rst-5e-12)/10e-6))'
+NRS='wn_rst/ceil((wn_rst-5e-12)/10e-6)<119.5e-9?(((14.4e-15+(wn_rst/ceil((wn_rst-5e-12)/10e-6))*50e-9)+floor((ceil((wn_rst-5e-12)/10e-6)-1)/2.0)*(14.4e-15+(wn_rst/ceil((wn_rst-5e-12)/10e-6))*100e-9))+(ceil((wn_rst-5e-12)/10e-6)/2-floor(ceil((wn_rst-5e-12)/10e-6)/2)==0?14.4e-15+(wn_rst/ceil((wn_rst-5e-12)/10e-6))*50e-9:0))/1:(((140e-9*(wn_rst/ceil((wn_rst-5e-12)/10e-6))+floor((ceil((wn_rst-5e-12)/10e-6)-1)/2.0)*(110e-9*(wn_rst/ceil((wn_rst-5e-12)/10e-6))))+(ceil((wn_rst-5e-12)/10e-6)/2-floor(ceil((wn_rst-5e-12)/10e-6)/2)==0?140e-9*(wn_rst/ceil((wn_rst-5e-12)/10e-6)):0))/1)/((((wn_rst/ceil((wn_rst-5e-12)/10e-6))*ceil((wn_rst-5e-12)/10e-6))*(wn_rst/ceil((wn_rst-5e-12)/10e-6)))*ceil((wn_rst-5e-12)/10e-6))' M=1

mnm4 x rst vss vss g45n1svt L=45e-9 W=wn_rst AD='wn_rst/ceil((wn_rst-5e-12)/10e-6)<119.5e-9?(floor(ceil((wn_rst-5e-12)/10e-6)/2.0)*(14.4e-15+(wn_rst/ceil((wn_rst-5e-12)/10e-6))*100e-9)+(ceil((wn_rst-5e-12)/10e-6)/2-floor(ceil((wn_rst-5e-12)/10e-6)/2)!=0?14.4e-15+(wn_rst/ceil((wn_rst-5e-12)/10e-6))*50e-9:0))/1:(floor(ceil((wn_rst-5e-12)/10e-6)/2.0)*(110e-9*(wn_rst/ceil((wn_rst-5e-12)/10e-6)))+(ceil((wn_rst-5e-12)/10e-6)/2-floor(ceil((wn_rst-5e-12)/10e-6)/2)!=0?140e-9*(wn_rst/ceil((wn_rst-5e-12)/10e-6)):0))/1'
+AS='wn_rst/ceil((wn_rst-5e-12)/10e-6)<119.5e-9?(((14.4e-15+(wn_rst/ceil((wn_rst-5e-12)/10e-6))*50e-9)+floor((ceil((wn_rst-5e-12)/10e-6)-1)/2.0)*(14.4e-15+(wn_rst/ceil((wn_rst-5e-12)/10e-6))*100e-9))+(ceil((wn_rst-5e-12)/10e-6)/2-floor(ceil((wn_rst-5e-12)/10e-6)/2)==0?14.4e-15+(wn_rst/ceil((wn_rst-5e-12)/10e-6))*50e-9:0))/1:((140e-9*(wn_rst/ceil((wn_rst-5e-12)/10e-6))+floor((ceil((wn_rst-5e-12)/10e-6)-1)/2.0)*(110e-9*(wn_rst/ceil((wn_rst-5e-12)/10e-6))))+(ceil((wn_rst-5e-12)/10e-6)/2-floor(ceil((wn_rst-5e-12)/10e-6)/2)==0?140e-9*(wn_rst/ceil((wn_rst-5e-12)/10e-6)):0))/1' PD='wn_rst/ceil((wn_rst-5e-12)/10e-6)<119.5e-9?(floor(ceil((wn_rst-5e-12)/10e-6)/2.0)*680e-9+(ceil((wn_rst-5e-12)/10e-6)/2-floor(ceil((wn_rst-5e-12)/10e-6)/2)!=0?580e-9:0))/1:(floor(ceil((wn_rst-5e-12)/10e-6)/2.0)*(220e-9+2*(wn_rst/ceil((wn_rst-5e-12)/10e-6)))+(ceil((wn_rst-5e-12)/10e-6)/2-floor(ceil((wn_rst-5e-12)/10e-6)/2)!=0?280e-9+2*(wn_rst/ceil((wn_rst-5e-12)/10e-6)):0))/1'
+PS='wn_rst/ceil((wn_rst-5e-12)/10e-6)<119.5e-9?((580e-9+floor((ceil((wn_rst-5e-12)/10e-6)-1)/2.0)*680e-9)+(ceil((wn_rst-5e-12)/10e-6)/2-floor(ceil((wn_rst-5e-12)/10e-6)/2)==0?580e-9:0))/1:(((280e-9+2*(wn_rst/ceil((wn_rst-5e-12)/10e-6)))+floor((ceil((wn_rst-5e-12)/10e-6)-1)/2.0)*(220e-9+2*(wn_rst/ceil((wn_rst-5e-12)/10e-6))))+(ceil((wn_rst-5e-12)/10e-6)/2-floor(ceil((wn_rst-5e-12)/10e-6)/2)==0?280e-9+2*(wn_rst/ceil((wn_rst-5e-12)/10e-6)):0))/1'
+NRD='wn_rst/ceil((wn_rst-5e-12)/10e-6)<119.5e-9?(floor(ceil((wn_rst-5e-12)/10e-6)/2.0)*(14.4e-15+(wn_rst/ceil((wn_rst-5e-12)/10e-6))*100e-9)+(ceil((wn_rst-5e-12)/10e-6)/2-floor(ceil((wn_rst-5e-12)/10e-6)/2)!=0?14.4e-15+(wn_rst/ceil((wn_rst-5e-12)/10e-6))*50e-9:0))/1:((floor(ceil((wn_rst-5e-12)/10e-6)/2.0)*(110e-9*(wn_rst/ceil((wn_rst-5e-12)/10e-6)))+(ceil((wn_rst-5e-12)/10e-6)/2-floor(ceil((wn_rst-5e-12)/10e-6)/2)!=0?140e-9*(wn_rst/ceil((wn_rst-5e-12)/10e-6)):0))/1)/((((wn_rst/ceil((wn_rst-5e-12)/10e-6))*ceil((wn_rst-5e-12)/10e-6))*(wn_rst/ceil((wn_rst-5e-12)/10e-6)))*ceil((wn_rst-5e-12)/10e-6))'
+NRS='wn_rst/ceil((wn_rst-5e-12)/10e-6)<119.5e-9?(((14.4e-15+(wn_rst/ceil((wn_rst-5e-12)/10e-6))*50e-9)+floor((ceil((wn_rst-5e-12)/10e-6)-1)/2.0)*(14.4e-15+(wn_rst/ceil((wn_rst-5e-12)/10e-6))*100e-9))+(ceil((wn_rst-5e-12)/10e-6)/2-floor(ceil((wn_rst-5e-12)/10e-6)/2)==0?14.4e-15+(wn_rst/ceil((wn_rst-5e-12)/10e-6))*50e-9:0))/1:(((140e-9*(wn_rst/ceil((wn_rst-5e-12)/10e-6))+floor((ceil((wn_rst-5e-12)/10e-6)-1)/2.0)*(110e-9*(wn_rst/ceil((wn_rst-5e-12)/10e-6))))+(ceil((wn_rst-5e-12)/10e-6)/2-floor(ceil((wn_rst-5e-12)/10e-6)/2)==0?140e-9*(wn_rst/ceil((wn_rst-5e-12)/10e-6)):0))/1)/((((wn_rst/ceil((wn_rst-5e-12)/10e-6))*ceil((wn_rst-5e-12)/10e-6))*(wn_rst/ceil((wn_rst-5e-12)/10e-6)))*ceil((wn_rst-5e-12)/10e-6))' M=1

mnm3 net21 x vss vss g45n1svt L=45e-9 W=wn_q AD='wn_q/ceil((wn_q-5e-12)/10e-6)<119.5e-9?(floor(ceil((wn_q-5e-12)/10e-6)/2.0)*(14.4e-15+(wn_q/ceil((wn_q-5e-12)/10e-6))*100e-9)+(ceil((wn_q-5e-12)/10e-6)/2-floor(ceil((wn_q-5e-12)/10e-6)/2)!=0?14.4e-15+(wn_q/ceil((wn_q-5e-12)/10e-6))*50e-9:0))/1:(floor(ceil((wn_q-5e-12)/10e-6)/2.0)*(110e-9*(wn_q/ceil((wn_q-5e-12)/10e-6)))+(ceil((wn_q-5e-12)/10e-6)/2-floor(ceil((wn_q-5e-12)/10e-6)/2)!=0?140e-9*(wn_q/ceil((wn_q-5e-12)/10e-6)):0))/1' AS='wn_q/ceil((wn_q-5e-12)/10e-6)<119.5e-9?(((14.4e-15+(wn_q/ceil((wn_q-5e-12)/10e-6))*50e-9)+floor((ceil((wn_q-5e-12)/10e-6)-1)/2.0)*(14.4e-15+(wn_q/ceil((wn_q-5e-12)/10e-6))*100e-9))+(ceil((wn_q-5e-12)/10e-6)/2-floor(ceil((wn_q-5e-12)/10e-6)/2)==0?14.4e-15+(wn_q/ceil((wn_q-5e-12)/10e-6))*50e-9:0))/1:((140e-9*(wn_q/ceil((wn_q-5e-12)/10e-6))+floor((ceil((wn_q-5e-12)/10e-6)-1)/2.0)*(110e-9*(wn_q/ceil((wn_q-5e-12)/10e-6))))+(ceil((wn_q-5e-12)/10e-6)/2-floor(ceil((wn_q-5e-12)/10e-6)/2)==0?140e-9*(wn_q/ceil((wn_q-5e-12)/10e-6)):0))/1'
+PD='wn_q/ceil((wn_q-5e-12)/10e-6)<119.5e-9?(floor(ceil((wn_q-5e-12)/10e-6)/2.0)*680e-9+(ceil((wn_q-5e-12)/10e-6)/2-floor(ceil((wn_q-5e-12)/10e-6)/2)!=0?580e-9:0))/1:(floor(ceil((wn_q-5e-12)/10e-6)/2.0)*(220e-9+2*(wn_q/ceil((wn_q-5e-12)/10e-6)))+(ceil((wn_q-5e-12)/10e-6)/2-floor(ceil((wn_q-5e-12)/10e-6)/2)!=0?280e-9+2*(wn_q/ceil((wn_q-5e-12)/10e-6)):0))/1' PS='wn_q/ceil((wn_q-5e-12)/10e-6)<119.5e-9?((580e-9+floor((ceil((wn_q-5e-12)/10e-6)-1)/2.0)*680e-9)+(ceil((wn_q-5e-12)/10e-6)/2-floor(ceil((wn_q-5e-12)/10e-6)/2)==0?580e-9:0))/1:(((280e-9+2*(wn_q/ceil((wn_q-5e-12)/10e-6)))+floor((ceil((wn_q-5e-12)/10e-6)-1)/2.0)*(220e-9+2*(wn_q/ceil((wn_q-5e-12)/10e-6))))+(ceil((wn_q-5e-12)/10e-6)/2-floor(ceil((wn_q-5e-12)/10e-6)/2)==0?280e-9+2*(wn_q/ceil((wn_q-5e-12)/10e-6)):0))/1'
+NRD='wn_q/ceil((wn_q-5e-12)/10e-6)<119.5e-9?(floor(ceil((wn_q-5e-12)/10e-6)/2.0)*(14.4e-15+(wn_q/ceil((wn_q-5e-12)/10e-6))*100e-9)+(ceil((wn_q-5e-12)/10e-6)/2-floor(ceil((wn_q-5e-12)/10e-6)/2)!=0?14.4e-15+(wn_q/ceil((wn_q-5e-12)/10e-6))*50e-9:0))/1:((floor(ceil((wn_q-5e-12)/10e-6)/2.0)*(110e-9*(wn_q/ceil((wn_q-5e-12)/10e-6)))+(ceil((wn_q-5e-12)/10e-6)/2-floor(ceil((wn_q-5e-12)/10e-6)/2)!=0?140e-9*(wn_q/ceil((wn_q-5e-12)/10e-6)):0))/1)/((((wn_q/ceil((wn_q-5e-12)/10e-6))*ceil((wn_q-5e-12)/10e-6))*(wn_q/ceil((wn_q-5e-12)/10e-6)))*ceil((wn_q-5e-12)/10e-6))'
+NRS='wn_q/ceil((wn_q-5e-12)/10e-6)<119.5e-9?(((14.4e-15+(wn_q/ceil((wn_q-5e-12)/10e-6))*50e-9)+floor((ceil((wn_q-5e-12)/10e-6)-1)/2.0)*(14.4e-15+(wn_q/ceil((wn_q-5e-12)/10e-6))*100e-9))+(ceil((wn_q-5e-12)/10e-6)/2-floor(ceil((wn_q-5e-12)/10e-6)/2)==0?14.4e-15+(wn_q/ceil((wn_q-5e-12)/10e-6))*50e-9:0))/1:(((140e-9*(wn_q/ceil((wn_q-5e-12)/10e-6))+floor((ceil((wn_q-5e-12)/10e-6)-1)/2.0)*(110e-9*(wn_q/ceil((wn_q-5e-12)/10e-6))))+(ceil((wn_q-5e-12)/10e-6)/2-floor(ceil((wn_q-5e-12)/10e-6)/2)==0?140e-9*(wn_q/ceil((wn_q-5e-12)/10e-6)):0))/1)/((((wn_q/ceil((wn_q-5e-12)/10e-6))*ceil((wn_q-5e-12)/10e-6))*(wn_q/ceil((wn_q-5e-12)/10e-6)))*ceil((wn_q-5e-12)/10e-6))' M=1

mnm2 q clk net21 vss g45n1svt L=45e-9 W=wn_clk AD='wn_clk/ceil((wn_clk-5e-12)/10e-6)<119.5e-9?(floor(ceil((wn_clk-5e-12)/10e-6)/2.0)*(14.4e-15+(wn_clk/ceil((wn_clk-5e-12)/10e-6))*100e-9)+(ceil((wn_clk-5e-12)/10e-6)/2-floor(ceil((wn_clk-5e-12)/10e-6)/2)!=0?14.4e-15+(wn_clk/ceil((wn_clk-5e-12)/10e-6))*50e-9:0))/1:(floor(ceil((wn_clk-5e-12)/10e-6)/2.0)*(110e-9*(wn_clk/ceil((wn_clk-5e-12)/10e-6)))+(ceil((wn_clk-5e-12)/10e-6)/2-floor(ceil((wn_clk-5e-12)/10e-6)/2)!=0?140e-9*(wn_clk/ceil((wn_clk-5e-12)/10e-6)):0))/1'
+AS='wn_clk/ceil((wn_clk-5e-12)/10e-6)<119.5e-9?(((14.4e-15+(wn_clk/ceil((wn_clk-5e-12)/10e-6))*50e-9)+floor((ceil((wn_clk-5e-12)/10e-6)-1)/2.0)*(14.4e-15+(wn_clk/ceil((wn_clk-5e-12)/10e-6))*100e-9))+(ceil((wn_clk-5e-12)/10e-6)/2-floor(ceil((wn_clk-5e-12)/10e-6)/2)==0?14.4e-15+(wn_clk/ceil((wn_clk-5e-12)/10e-6))*50e-9:0))/1:((140e-9*(wn_clk/ceil((wn_clk-5e-12)/10e-6))+floor((ceil((wn_clk-5e-12)/10e-6)-1)/2.0)*(110e-9*(wn_clk/ceil((wn_clk-5e-12)/10e-6))))+(ceil((wn_clk-5e-12)/10e-6)/2-floor(ceil((wn_clk-5e-12)/10e-6)/2)==0?140e-9*(wn_clk/ceil((wn_clk-5e-12)/10e-6)):0))/1' PD='wn_clk/ceil((wn_clk-5e-12)/10e-6)<119.5e-9?(floor(ceil((wn_clk-5e-12)/10e-6)/2.0)*680e-9+(ceil((wn_clk-5e-12)/10e-6)/2-floor(ceil((wn_clk-5e-12)/10e-6)/2)!=0?580e-9:0))/1:(floor(ceil((wn_clk-5e-12)/10e-6)/2.0)*(220e-9+2*(wn_clk/ceil((wn_clk-5e-12)/10e-6)))+(ceil((wn_clk-5e-12)/10e-6)/2-floor(ceil((wn_clk-5e-12)/10e-6)/2)!=0?280e-9+2*(wn_clk/ceil((wn_clk-5e-12)/10e-6)):0))/1'
+PS='wn_clk/ceil((wn_clk-5e-12)/10e-6)<119.5e-9?((580e-9+floor((ceil((wn_clk-5e-12)/10e-6)-1)/2.0)*680e-9)+(ceil((wn_clk-5e-12)/10e-6)/2-floor(ceil((wn_clk-5e-12)/10e-6)/2)==0?580e-9:0))/1:(((280e-9+2*(wn_clk/ceil((wn_clk-5e-12)/10e-6)))+floor((ceil((wn_clk-5e-12)/10e-6)-1)/2.0)*(220e-9+2*(wn_clk/ceil((wn_clk-5e-12)/10e-6))))+(ceil((wn_clk-5e-12)/10e-6)/2-floor(ceil((wn_clk-5e-12)/10e-6)/2)==0?280e-9+2*(wn_clk/ceil((wn_clk-5e-12)/10e-6)):0))/1'
+NRD='wn_clk/ceil((wn_clk-5e-12)/10e-6)<119.5e-9?(floor(ceil((wn_clk-5e-12)/10e-6)/2.0)*(14.4e-15+(wn_clk/ceil((wn_clk-5e-12)/10e-6))*100e-9)+(ceil((wn_clk-5e-12)/10e-6)/2-floor(ceil((wn_clk-5e-12)/10e-6)/2)!=0?14.4e-15+(wn_clk/ceil((wn_clk-5e-12)/10e-6))*50e-9:0))/1:((floor(ceil((wn_clk-5e-12)/10e-6)/2.0)*(110e-9*(wn_clk/ceil((wn_clk-5e-12)/10e-6)))+(ceil((wn_clk-5e-12)/10e-6)/2-floor(ceil((wn_clk-5e-12)/10e-6)/2)!=0?140e-9*(wn_clk/ceil((wn_clk-5e-12)/10e-6)):0))/1)/((((wn_clk/ceil((wn_clk-5e-12)/10e-6))*ceil((wn_clk-5e-12)/10e-6))*(wn_clk/ceil((wn_clk-5e-12)/10e-6)))*ceil((wn_clk-5e-12)/10e-6))'
+NRS='wn_clk/ceil((wn_clk-5e-12)/10e-6)<119.5e-9?(((14.4e-15+(wn_clk/ceil((wn_clk-5e-12)/10e-6))*50e-9)+floor((ceil((wn_clk-5e-12)/10e-6)-1)/2.0)*(14.4e-15+(wn_clk/ceil((wn_clk-5e-12)/10e-6))*100e-9))+(ceil((wn_clk-5e-12)/10e-6)/2-floor(ceil((wn_clk-5e-12)/10e-6)/2)==0?14.4e-15+(wn_clk/ceil((wn_clk-5e-12)/10e-6))*50e-9:0))/1:(((140e-9*(wn_clk/ceil((wn_clk-5e-12)/10e-6))+floor((ceil((wn_clk-5e-12)/10e-6)-1)/2.0)*(110e-9*(wn_clk/ceil((wn_clk-5e-12)/10e-6))))+(ceil((wn_clk-5e-12)/10e-6)/2-floor(ceil((wn_clk-5e-12)/10e-6)/2)==0?140e-9*(wn_clk/ceil((wn_clk-5e-12)/10e-6)):0))/1)/((((wn_clk/ceil((wn_clk-5e-12)/10e-6))*ceil((wn_clk-5e-12)/10e-6))*(wn_clk/ceil((wn_clk-5e-12)/10e-6)))*ceil((wn_clk-5e-12)/10e-6))' M=1

mnm1 net9 d vss vss g45n1svt L=45e-9 W=wn_d AD='wn_d/ceil((wn_d-5e-12)/10e-6)<119.5e-9?(floor(ceil((wn_d-5e-12)/10e-6)/2.0)*(14.4e-15+(wn_d/ceil((wn_d-5e-12)/10e-6))*100e-9)+(ceil((wn_d-5e-12)/10e-6)/2-floor(ceil((wn_d-5e-12)/10e-6)/2)!=0?14.4e-15+(wn_d/ceil((wn_d-5e-12)/10e-6))*50e-9:0))/1:(floor(ceil((wn_d-5e-12)/10e-6)/2.0)*(110e-9*(wn_d/ceil((wn_d-5e-12)/10e-6)))+(ceil((wn_d-5e-12)/10e-6)/2-floor(ceil((wn_d-5e-12)/10e-6)/2)!=0?140e-9*(wn_d/ceil((wn_d-5e-12)/10e-6)):0))/1'
+AS='wn_d/ceil((wn_d-5e-12)/10e-6)<119.5e-9?(((14.4e-15+(wn_d/ceil((wn_d-5e-12)/10e-6))*50e-9)+floor((ceil((wn_d-5e-12)/10e-6)-1)/2.0)*(14.4e-15+(wn_d/ceil((wn_d-5e-12)/10e-6))*100e-9))+(ceil((wn_d-5e-12)/10e-6)/2-floor(ceil((wn_d-5e-12)/10e-6)/2)==0?14.4e-15+(wn_d/ceil((wn_d-5e-12)/10e-6))*50e-9:0))/1:((140e-9*(wn_d/ceil((wn_d-5e-12)/10e-6))+floor((ceil((wn_d-5e-12)/10e-6)-1)/2.0)*(110e-9*(wn_d/ceil((wn_d-5e-12)/10e-6))))+(ceil((wn_d-5e-12)/10e-6)/2-floor(ceil((wn_d-5e-12)/10e-6)/2)==0?140e-9*(wn_d/ceil((wn_d-5e-12)/10e-6)):0))/1' PD='wn_d/ceil((wn_d-5e-12)/10e-6)<119.5e-9?(floor(ceil((wn_d-5e-12)/10e-6)/2.0)*680e-9+(ceil((wn_d-5e-12)/10e-6)/2-floor(ceil((wn_d-5e-12)/10e-6)/2)!=0?580e-9:0))/1:(floor(ceil((wn_d-5e-12)/10e-6)/2.0)*(220e-9+2*(wn_d/ceil((wn_d-5e-12)/10e-6)))+(ceil((wn_d-5e-12)/10e-6)/2-floor(ceil((wn_d-5e-12)/10e-6)/2)!=0?280e-9+2*(wn_d/ceil((wn_d-5e-12)/10e-6)):0))/1'
+PS='wn_d/ceil((wn_d-5e-12)/10e-6)<119.5e-9?((580e-9+floor((ceil((wn_d-5e-12)/10e-6)-1)/2.0)*680e-9)+(ceil((wn_d-5e-12)/10e-6)/2-floor(ceil((wn_d-5e-12)/10e-6)/2)==0?580e-9:0))/1:(((280e-9+2*(wn_d/ceil((wn_d-5e-12)/10e-6)))+floor((ceil((wn_d-5e-12)/10e-6)-1)/2.0)*(220e-9+2*(wn_d/ceil((wn_d-5e-12)/10e-6))))+(ceil((wn_d-5e-12)/10e-6)/2-floor(ceil((wn_d-5e-12)/10e-6)/2)==0?280e-9+2*(wn_d/ceil((wn_d-5e-12)/10e-6)):0))/1'
+NRD='wn_d/ceil((wn_d-5e-12)/10e-6)<119.5e-9?(floor(ceil((wn_d-5e-12)/10e-6)/2.0)*(14.4e-15+(wn_d/ceil((wn_d-5e-12)/10e-6))*100e-9)+(ceil((wn_d-5e-12)/10e-6)/2-floor(ceil((wn_d-5e-12)/10e-6)/2)!=0?14.4e-15+(wn_d/ceil((wn_d-5e-12)/10e-6))*50e-9:0))/1:((floor(ceil((wn_d-5e-12)/10e-6)/2.0)*(110e-9*(wn_d/ceil((wn_d-5e-12)/10e-6)))+(ceil((wn_d-5e-12)/10e-6)/2-floor(ceil((wn_d-5e-12)/10e-6)/2)!=0?140e-9*(wn_d/ceil((wn_d-5e-12)/10e-6)):0))/1)/((((wn_d/ceil((wn_d-5e-12)/10e-6))*ceil((wn_d-5e-12)/10e-6))*(wn_d/ceil((wn_d-5e-12)/10e-6)))*ceil((wn_d-5e-12)/10e-6))'
+NRS='wn_d/ceil((wn_d-5e-12)/10e-6)<119.5e-9?(((14.4e-15+(wn_d/ceil((wn_d-5e-12)/10e-6))*50e-9)+floor((ceil((wn_d-5e-12)/10e-6)-1)/2.0)*(14.4e-15+(wn_d/ceil((wn_d-5e-12)/10e-6))*100e-9))+(ceil((wn_d-5e-12)/10e-6)/2-floor(ceil((wn_d-5e-12)/10e-6)/2)==0?14.4e-15+(wn_d/ceil((wn_d-5e-12)/10e-6))*50e-9:0))/1:(((140e-9*(wn_d/ceil((wn_d-5e-12)/10e-6))+floor((ceil((wn_d-5e-12)/10e-6)-1)/2.0)*(110e-9*(wn_d/ceil((wn_d-5e-12)/10e-6))))+(ceil((wn_d-5e-12)/10e-6)/2-floor(ceil((wn_d-5e-12)/10e-6)/2)==0?140e-9*(wn_d/ceil((wn_d-5e-12)/10e-6)):0))/1)/((((wn_d/ceil((wn_d-5e-12)/10e-6))*ceil((wn_d-5e-12)/10e-6))*(wn_d/ceil((wn_d-5e-12)/10e-6)))*ceil((wn_d-5e-12)/10e-6))' M=1

mnm0 x clk_bar net9 vss g45n1svt L=45e-9 W=wn_clk AD='wn_clk/ceil((wn_clk-5e-12)/10e-6)<119.5e-9?(floor(ceil((wn_clk-5e-12)/10e-6)/2.0)*(14.4e-15+(wn_clk/ceil((wn_clk-5e-12)/10e-6))*100e-9)+(ceil((wn_clk-5e-12)/10e-6)/2-floor(ceil((wn_clk-5e-12)/10e-6)/2)!=0?14.4e-15+(wn_clk/ceil((wn_clk-5e-12)/10e-6))*50e-9:0))/1:(floor(ceil((wn_clk-5e-12)/10e-6)/2.0)*(110e-9*(wn_clk/ceil((wn_clk-5e-12)/10e-6)))+(ceil((wn_clk-5e-12)/10e-6)/2-floor(ceil((wn_clk-5e-12)/10e-6)/2)!=0?140e-9*(wn_clk/ceil((wn_clk-5e-12)/10e-6)):0))/1'
+AS='wn_clk/ceil((wn_clk-5e-12)/10e-6)<119.5e-9?(((14.4e-15+(wn_clk/ceil((wn_clk-5e-12)/10e-6))*50e-9)+floor((ceil((wn_clk-5e-12)/10e-6)-1)/2.0)*(14.4e-15+(wn_clk/ceil((wn_clk-5e-12)/10e-6))*100e-9))+(ceil((wn_clk-5e-12)/10e-6)/2-floor(ceil((wn_clk-5e-12)/10e-6)/2)==0?14.4e-15+(wn_clk/ceil((wn_clk-5e-12)/10e-6))*50e-9:0))/1:((140e-9*(wn_clk/ceil((wn_clk-5e-12)/10e-6))+floor((ceil((wn_clk-5e-12)/10e-6)-1)/2.0)*(110e-9*(wn_clk/ceil((wn_clk-5e-12)/10e-6))))+(ceil((wn_clk-5e-12)/10e-6)/2-floor(ceil((wn_clk-5e-12)/10e-6)/2)==0?140e-9*(wn_clk/ceil((wn_clk-5e-12)/10e-6)):0))/1' PD='wn_clk/ceil((wn_clk-5e-12)/10e-6)<119.5e-9?(floor(ceil((wn_clk-5e-12)/10e-6)/2.0)*680e-9+(ceil((wn_clk-5e-12)/10e-6)/2-floor(ceil((wn_clk-5e-12)/10e-6)/2)!=0?580e-9:0))/1:(floor(ceil((wn_clk-5e-12)/10e-6)/2.0)*(220e-9+2*(wn_clk/ceil((wn_clk-5e-12)/10e-6)))+(ceil((wn_clk-5e-12)/10e-6)/2-floor(ceil((wn_clk-5e-12)/10e-6)/2)!=0?280e-9+2*(wn_clk/ceil((wn_clk-5e-12)/10e-6)):0))/1'
+PS='wn_clk/ceil((wn_clk-5e-12)/10e-6)<119.5e-9?((580e-9+floor((ceil((wn_clk-5e-12)/10e-6)-1)/2.0)*680e-9)+(ceil((wn_clk-5e-12)/10e-6)/2-floor(ceil((wn_clk-5e-12)/10e-6)/2)==0?580e-9:0))/1:(((280e-9+2*(wn_clk/ceil((wn_clk-5e-12)/10e-6)))+floor((ceil((wn_clk-5e-12)/10e-6)-1)/2.0)*(220e-9+2*(wn_clk/ceil((wn_clk-5e-12)/10e-6))))+(ceil((wn_clk-5e-12)/10e-6)/2-floor(ceil((wn_clk-5e-12)/10e-6)/2)==0?280e-9+2*(wn_clk/ceil((wn_clk-5e-12)/10e-6)):0))/1'
+NRD='wn_clk/ceil((wn_clk-5e-12)/10e-6)<119.5e-9?(floor(ceil((wn_clk-5e-12)/10e-6)/2.0)*(14.4e-15+(wn_clk/ceil((wn_clk-5e-12)/10e-6))*100e-9)+(ceil((wn_clk-5e-12)/10e-6)/2-floor(ceil((wn_clk-5e-12)/10e-6)/2)!=0?14.4e-15+(wn_clk/ceil((wn_clk-5e-12)/10e-6))*50e-9:0))/1:((floor(ceil((wn_clk-5e-12)/10e-6)/2.0)*(110e-9*(wn_clk/ceil((wn_clk-5e-12)/10e-6)))+(ceil((wn_clk-5e-12)/10e-6)/2-floor(ceil((wn_clk-5e-12)/10e-6)/2)!=0?140e-9*(wn_clk/ceil((wn_clk-5e-12)/10e-6)):0))/1)/((((wn_clk/ceil((wn_clk-5e-12)/10e-6))*ceil((wn_clk-5e-12)/10e-6))*(wn_clk/ceil((wn_clk-5e-12)/10e-6)))*ceil((wn_clk-5e-12)/10e-6))'
+NRS='wn_clk/ceil((wn_clk-5e-12)/10e-6)<119.5e-9?(((14.4e-15+(wn_clk/ceil((wn_clk-5e-12)/10e-6))*50e-9)+floor((ceil((wn_clk-5e-12)/10e-6)-1)/2.0)*(14.4e-15+(wn_clk/ceil((wn_clk-5e-12)/10e-6))*100e-9))+(ceil((wn_clk-5e-12)/10e-6)/2-floor(ceil((wn_clk-5e-12)/10e-6)/2)==0?14.4e-15+(wn_clk/ceil((wn_clk-5e-12)/10e-6))*50e-9:0))/1:(((140e-9*(wn_clk/ceil((wn_clk-5e-12)/10e-6))+floor((ceil((wn_clk-5e-12)/10e-6)-1)/2.0)*(110e-9*(wn_clk/ceil((wn_clk-5e-12)/10e-6))))+(ceil((wn_clk-5e-12)/10e-6)/2-floor(ceil((wn_clk-5e-12)/10e-6)/2)==0?140e-9*(wn_clk/ceil((wn_clk-5e-12)/10e-6)):0))/1)/((((wn_clk/ceil((wn_clk-5e-12)/10e-6))*ceil((wn_clk-5e-12)/10e-6))*(wn_clk/ceil((wn_clk-5e-12)/10e-6)))*ceil((wn_clk-5e-12)/10e-6))' M=1

Cq  q  vss  10f
Cx  x  vss  10f

* ----------------------------------------------------------
* TRANSIENT ANALYSIS + MEASURES
* ----------------------------------------------------------
.tran 1p 40n

* Basic probes
.probe v(d) v(clk) v(clk_bar) v(rst) v(x) v(q)

* Simple timing measures (example: Q rising delay from D)
.measure tran t_d_rise  trig v(d)  val=0.55 rise=1
+                        targ v(q)  val=0.55 rise=1

.measure tran t_d_fall  trig v(d)  val=0.55 fall=1
+                        targ v(q)  val=0.55 fall=1

.END
