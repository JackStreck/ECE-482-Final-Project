* resm11_pcell_1.sp
.subckt resm11_pcell_1 P N
R1 P N 3.5m
.ends resm11_pcell_1

.subckt resm11_pcell_01 P N
R1 P N 3.5m
.ends resm11_pcell_01

.subckt resm11_pcell_0 P N
R1 P N 3.5m
.ends resm11_pcell_0

