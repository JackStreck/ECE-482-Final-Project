ECE 482 PROJECT TESTBENCH
.lib '/class/ece482/gpdk045_mos' SS
.include "resm11_pcell_1.sp"

*The following parameter can be modified.
.param nom_vdd = 1.1

*The following parameters cannot be modified.
.param tstart = 1n
.param TCK = 4n
.param trf_ck = 200p
.param trf_ip_reset = 200p
.param reset_pw = 6n
.param CK_pw = 0.5*TCK
.param reset_delay = 1n
.param reset_delay2 = 10n
.param sim_end = 11*TCK
.param input_delay = 9.5n
.param input_delay2 = 9.7n
.param input_delay3 = 9.2n
.param input_delay4 = 9.8n
.param input_pw = 1*TCK
.param offset_ip = 1n

*Put your extracted netlist below this comment

** Library name: test2
** Cell name: level_shifter_1_1_to_1_8
** View name: schematic
.subckt level_shifter_1_1_to_1_8 bio bio_bar b_core b_core_bar vdd vss
m1 bio b_core_bar vss vss g45n2svt L=150e-9 W=640e-9 AD='640e-9/ceil(63.9995e-3)<119.5e-9?(floor(ceil(63.9995e-3)/2.0)*(14.4e-15+(640e-9/ceil(63.9995e-3))*100e-9)+(ceil(63.9995e-3)/2-floor(ceil(63.9995e-3)/2)!=0?14.4e-15+(640e-9/ceil(63.9995e-3))*50e-9:0))/1:(floor(ceil(63.9995e-3)/2.0)*(200e-9*(640e-9/ceil(63.9995e-3)))+(ceil(63.9995e-3)/2-floor(ceil(63.9995e-3)/2)!=0?150e-9*(640e-9/ceil(63.9995e-3)):0))/1' AS='640e-9/ceil(63.9995e-3)<119.5e-9?(((14.4e-15+(640e-9/ceil(63.9995e-3))*50e-9)+floor((ceil(63.9995e-3)-1)/2.0)*(14.4e-15+(640e-9/ceil(63.9995e-3))*100e-9))+(ceil(63.9995e-3)/2-floor(ceil(63.9995e-3)/2)==0?14.4e-15+(640e-9/ceil(63.9995e-3))*50e-9:0))/1:((150e-9*(640e-9/ceil(63.9995e-3))+floor((ceil(63.9995e-3)-1)/2.0)*(200e-9*(640e-9/ceil(63.9995e-3))))+(ceil(63.9995e-3)/2-floor(ceil(63.9995e-3)/2)==0?150e-9*(640e-9/ceil(63.9995e-3)):0))/1'
+PD='640e-9/ceil(63.9995e-3)<119.5e-9?(floor(ceil(63.9995e-3)/2.0)*680e-9+(ceil(63.9995e-3)/2-floor(ceil(63.9995e-3)/2)!=0?580e-9:0))/1:(floor(ceil(63.9995e-3)/2.0)*(400e-9+2*(640e-9/ceil(63.9995e-3)))+(ceil(63.9995e-3)/2-floor(ceil(63.9995e-3)/2)!=0?300e-9+2*(640e-9/ceil(63.9995e-3)):0))/1' PS='640e-9/ceil(63.9995e-3)<119.5e-9?((580e-9+floor((ceil(63.9995e-3)-1)/2.0)*680e-9)+(ceil(63.9995e-3)/2-floor(ceil(63.9995e-3)/2)==0?580e-9:0))/1:(((300e-9+2*(640e-9/ceil(63.9995e-3)))+floor((ceil(63.9995e-3)-1)/2.0)*(400e-9+2*(640e-9/ceil(63.9995e-3))))+(ceil(63.9995e-3)/2-floor(ceil(63.9995e-3)/2)==0?300e-9+2*(640e-9/ceil(63.9995e-3)):0))/1'
+NRD='640e-9/ceil(63.9995e-3)<119.5e-9?(floor(ceil(63.9995e-3)/2.0)*(14.4e-15+(640e-9/ceil(63.9995e-3))*100e-9)+(ceil(63.9995e-3)/2-floor(ceil(63.9995e-3)/2)!=0?14.4e-15+(640e-9/ceil(63.9995e-3))*50e-9:0))/1:((floor(ceil(63.9995e-3)/2.0)*(200e-9*(640e-9/ceil(63.9995e-3)))+(ceil(63.9995e-3)/2-floor(ceil(63.9995e-3)/2)!=0?150e-9*(640e-9/ceil(63.9995e-3)):0))/1)/((((640e-9/ceil(63.9995e-3))*ceil(63.9995e-3))*(640e-9/ceil(63.9995e-3)))*ceil(63.9995e-3))' NRS='640e-9/ceil(63.9995e-3)<119.5e-9?(((14.4e-15+(640e-9/ceil(63.9995e-3))*50e-9)+floor((ceil(63.9995e-3)-1)/2.0)*(14.4e-15+(640e-9/ceil(63.9995e-3))*100e-9))+(ceil(63.9995e-3)/2-floor(ceil(63.9995e-3)/2)==0?14.4e-15+(640e-9/ceil(63.9995e-3))*50e-9:0))/1:(((150e-9*(640e-9/ceil(63.9995e-3))+floor((ceil(63.9995e-3)-1)/2.0)*(200e-9*(640e-9/ceil(63.9995e-3))))+(ceil(63.9995e-3)/2-floor(ceil(63.9995e-3)/2)==0?150e-9*(640e-9/ceil(63.9995e-3)):0))/1)/((((640e-9/ceil(63.9995e-3))*ceil(63.9995e-3))*(640e-9/ceil(63.9995e-3)))*ceil(63.9995e-3))' M=1
m0 bio_bar b_core vss vss g45n2svt L=150e-9 W=640e-9 AD='640e-9/ceil(63.9995e-3)<119.5e-9?(floor(ceil(63.9995e-3)/2.0)*(14.4e-15+(640e-9/ceil(63.9995e-3))*100e-9)+(ceil(63.9995e-3)/2-floor(ceil(63.9995e-3)/2)!=0?14.4e-15+(640e-9/ceil(63.9995e-3))*50e-9:0))/1:(floor(ceil(63.9995e-3)/2.0)*(200e-9*(640e-9/ceil(63.9995e-3)))+(ceil(63.9995e-3)/2-floor(ceil(63.9995e-3)/2)!=0?150e-9*(640e-9/ceil(63.9995e-3)):0))/1' AS='640e-9/ceil(63.9995e-3)<119.5e-9?(((14.4e-15+(640e-9/ceil(63.9995e-3))*50e-9)+floor((ceil(63.9995e-3)-1)/2.0)*(14.4e-15+(640e-9/ceil(63.9995e-3))*100e-9))+(ceil(63.9995e-3)/2-floor(ceil(63.9995e-3)/2)==0?14.4e-15+(640e-9/ceil(63.9995e-3))*50e-9:0))/1:((150e-9*(640e-9/ceil(63.9995e-3))+floor((ceil(63.9995e-3)-1)/2.0)*(200e-9*(640e-9/ceil(63.9995e-3))))+(ceil(63.9995e-3)/2-floor(ceil(63.9995e-3)/2)==0?150e-9*(640e-9/ceil(63.9995e-3)):0))/1'
+PD='640e-9/ceil(63.9995e-3)<119.5e-9?(floor(ceil(63.9995e-3)/2.0)*680e-9+(ceil(63.9995e-3)/2-floor(ceil(63.9995e-3)/2)!=0?580e-9:0))/1:(floor(ceil(63.9995e-3)/2.0)*(400e-9+2*(640e-9/ceil(63.9995e-3)))+(ceil(63.9995e-3)/2-floor(ceil(63.9995e-3)/2)!=0?300e-9+2*(640e-9/ceil(63.9995e-3)):0))/1' PS='640e-9/ceil(63.9995e-3)<119.5e-9?((580e-9+floor((ceil(63.9995e-3)-1)/2.0)*680e-9)+(ceil(63.9995e-3)/2-floor(ceil(63.9995e-3)/2)==0?580e-9:0))/1:(((300e-9+2*(640e-9/ceil(63.9995e-3)))+floor((ceil(63.9995e-3)-1)/2.0)*(400e-9+2*(640e-9/ceil(63.9995e-3))))+(ceil(63.9995e-3)/2-floor(ceil(63.9995e-3)/2)==0?300e-9+2*(640e-9/ceil(63.9995e-3)):0))/1'
+NRD='640e-9/ceil(63.9995e-3)<119.5e-9?(floor(ceil(63.9995e-3)/2.0)*(14.4e-15+(640e-9/ceil(63.9995e-3))*100e-9)+(ceil(63.9995e-3)/2-floor(ceil(63.9995e-3)/2)!=0?14.4e-15+(640e-9/ceil(63.9995e-3))*50e-9:0))/1:((floor(ceil(63.9995e-3)/2.0)*(200e-9*(640e-9/ceil(63.9995e-3)))+(ceil(63.9995e-3)/2-floor(ceil(63.9995e-3)/2)!=0?150e-9*(640e-9/ceil(63.9995e-3)):0))/1)/((((640e-9/ceil(63.9995e-3))*ceil(63.9995e-3))*(640e-9/ceil(63.9995e-3)))*ceil(63.9995e-3))' NRS='640e-9/ceil(63.9995e-3)<119.5e-9?(((14.4e-15+(640e-9/ceil(63.9995e-3))*50e-9)+floor((ceil(63.9995e-3)-1)/2.0)*(14.4e-15+(640e-9/ceil(63.9995e-3))*100e-9))+(ceil(63.9995e-3)/2-floor(ceil(63.9995e-3)/2)==0?14.4e-15+(640e-9/ceil(63.9995e-3))*50e-9:0))/1:(((150e-9*(640e-9/ceil(63.9995e-3))+floor((ceil(63.9995e-3)-1)/2.0)*(200e-9*(640e-9/ceil(63.9995e-3))))+(ceil(63.9995e-3)/2-floor(ceil(63.9995e-3)/2)==0?150e-9*(640e-9/ceil(63.9995e-3)):0))/1)/((((640e-9/ceil(63.9995e-3))*ceil(63.9995e-3))*(640e-9/ceil(63.9995e-3)))*ceil(63.9995e-3))' M=1
mpm1 bio bio_bar vdd vdd g45p2svt L=150e-9 W=480e-9 AD='480e-9/ceil(47.9995e-3)<119.5e-9?(floor(ceil(47.9995e-3)/2.0)*(14.4e-15+(480e-9/ceil(47.9995e-3))*100e-9)+(ceil(47.9995e-3)/2-floor(ceil(47.9995e-3)/2)!=0?14.4e-15+(480e-9/ceil(47.9995e-3))*50e-9:0))/1:(floor(ceil(47.9995e-3)/2.0)*(110e-9*(480e-9/ceil(47.9995e-3)))+(ceil(47.9995e-3)/2-floor(ceil(47.9995e-3)/2)!=0?140e-9*(480e-9/ceil(47.9995e-3)):0))/1' AS='480e-9/ceil(47.9995e-3)<119.5e-9?(((14.4e-15+(480e-9/ceil(47.9995e-3))*50e-9)+floor((ceil(47.9995e-3)-1)/2.0)*(14.4e-15+(480e-9/ceil(47.9995e-3))*100e-9))+(ceil(47.9995e-3)/2-floor(ceil(47.9995e-3)/2)==0?14.4e-15+(480e-9/ceil(47.9995e-3))*50e-9:0))/1:((140e-9*(480e-9/ceil(47.9995e-3))+floor((ceil(47.9995e-3)-1)/2.0)*(110e-9*(480e-9/ceil(47.9995e-3))))+(ceil(47.9995e-3)/2-floor(ceil(47.9995e-3)/2)==0?140e-9*(480e-9/ceil(47.9995e-3)):0))/1'
+PD='480e-9/ceil(47.9995e-3)<119.5e-9?(floor(ceil(47.9995e-3)/2.0)*680e-9+(ceil(47.9995e-3)/2-floor(ceil(47.9995e-3)/2)!=0?580e-9:0))/1:(floor(ceil(47.9995e-3)/2.0)*(220e-9+2*(480e-9/ceil(47.9995e-3)))+(ceil(47.9995e-3)/2-floor(ceil(47.9995e-3)/2)!=0?280e-9+2*(480e-9/ceil(47.9995e-3)):0))/1' PS='480e-9/ceil(47.9995e-3)<119.5e-9?((580e-9+floor((ceil(47.9995e-3)-1)/2.0)*680e-9)+(ceil(47.9995e-3)/2-floor(ceil(47.9995e-3)/2)==0?580e-9:0))/1:(((280e-9+2*(480e-9/ceil(47.9995e-3)))+floor((ceil(47.9995e-3)-1)/2.0)*(220e-9+2*(480e-9/ceil(47.9995e-3))))+(ceil(47.9995e-3)/2-floor(ceil(47.9995e-3)/2)==0?280e-9+2*(480e-9/ceil(47.9995e-3)):0))/1'
+NRD='480e-9/ceil(47.9995e-3)<119.5e-9?(floor(ceil(47.9995e-3)/2.0)*(14.4e-15+(480e-9/ceil(47.9995e-3))*100e-9)+(ceil(47.9995e-3)/2-floor(ceil(47.9995e-3)/2)!=0?14.4e-15+(480e-9/ceil(47.9995e-3))*50e-9:0))/1:((floor(ceil(47.9995e-3)/2.0)*(110e-9*(480e-9/ceil(47.9995e-3)))+(ceil(47.9995e-3)/2-floor(ceil(47.9995e-3)/2)!=0?140e-9*(480e-9/ceil(47.9995e-3)):0))/1)/((((480e-9/ceil(47.9995e-3))*ceil(47.9995e-3))*(480e-9/ceil(47.9995e-3)))*ceil(47.9995e-3))' NRS='480e-9/ceil(47.9995e-3)<119.5e-9?(((14.4e-15+(480e-9/ceil(47.9995e-3))*50e-9)+floor((ceil(47.9995e-3)-1)/2.0)*(14.4e-15+(480e-9/ceil(47.9995e-3))*100e-9))+(ceil(47.9995e-3)/2-floor(ceil(47.9995e-3)/2)==0?14.4e-15+(480e-9/ceil(47.9995e-3))*50e-9:0))/1:(((140e-9*(480e-9/ceil(47.9995e-3))+floor((ceil(47.9995e-3)-1)/2.0)*(110e-9*(480e-9/ceil(47.9995e-3))))+(ceil(47.9995e-3)/2-floor(ceil(47.9995e-3)/2)==0?140e-9*(480e-9/ceil(47.9995e-3)):0))/1)/((((480e-9/ceil(47.9995e-3))*ceil(47.9995e-3))*(480e-9/ceil(47.9995e-3)))*ceil(47.9995e-3))' M=1
mpm0 bio_bar bio vdd vdd g45p2svt L=150e-9 W=480e-9 AD='480e-9/ceil(47.9995e-3)<119.5e-9?(floor(ceil(47.9995e-3)/2.0)*(14.4e-15+(480e-9/ceil(47.9995e-3))*100e-9)+(ceil(47.9995e-3)/2-floor(ceil(47.9995e-3)/2)!=0?14.4e-15+(480e-9/ceil(47.9995e-3))*50e-9:0))/1:(floor(ceil(47.9995e-3)/2.0)*(110e-9*(480e-9/ceil(47.9995e-3)))+(ceil(47.9995e-3)/2-floor(ceil(47.9995e-3)/2)!=0?140e-9*(480e-9/ceil(47.9995e-3)):0))/1' AS='480e-9/ceil(47.9995e-3)<119.5e-9?(((14.4e-15+(480e-9/ceil(47.9995e-3))*50e-9)+floor((ceil(47.9995e-3)-1)/2.0)*(14.4e-15+(480e-9/ceil(47.9995e-3))*100e-9))+(ceil(47.9995e-3)/2-floor(ceil(47.9995e-3)/2)==0?14.4e-15+(480e-9/ceil(47.9995e-3))*50e-9:0))/1:((140e-9*(480e-9/ceil(47.9995e-3))+floor((ceil(47.9995e-3)-1)/2.0)*(110e-9*(480e-9/ceil(47.9995e-3))))+(ceil(47.9995e-3)/2-floor(ceil(47.9995e-3)/2)==0?140e-9*(480e-9/ceil(47.9995e-3)):0))/1'
+PD='480e-9/ceil(47.9995e-3)<119.5e-9?(floor(ceil(47.9995e-3)/2.0)*680e-9+(ceil(47.9995e-3)/2-floor(ceil(47.9995e-3)/2)!=0?580e-9:0))/1:(floor(ceil(47.9995e-3)/2.0)*(220e-9+2*(480e-9/ceil(47.9995e-3)))+(ceil(47.9995e-3)/2-floor(ceil(47.9995e-3)/2)!=0?280e-9+2*(480e-9/ceil(47.9995e-3)):0))/1' PS='480e-9/ceil(47.9995e-3)<119.5e-9?((580e-9+floor((ceil(47.9995e-3)-1)/2.0)*680e-9)+(ceil(47.9995e-3)/2-floor(ceil(47.9995e-3)/2)==0?580e-9:0))/1:(((280e-9+2*(480e-9/ceil(47.9995e-3)))+floor((ceil(47.9995e-3)-1)/2.0)*(220e-9+2*(480e-9/ceil(47.9995e-3))))+(ceil(47.9995e-3)/2-floor(ceil(47.9995e-3)/2)==0?280e-9+2*(480e-9/ceil(47.9995e-3)):0))/1'
+NRD='480e-9/ceil(47.9995e-3)<119.5e-9?(floor(ceil(47.9995e-3)/2.0)*(14.4e-15+(480e-9/ceil(47.9995e-3))*100e-9)+(ceil(47.9995e-3)/2-floor(ceil(47.9995e-3)/2)!=0?14.4e-15+(480e-9/ceil(47.9995e-3))*50e-9:0))/1:((floor(ceil(47.9995e-3)/2.0)*(110e-9*(480e-9/ceil(47.9995e-3)))+(ceil(47.9995e-3)/2-floor(ceil(47.9995e-3)/2)!=0?140e-9*(480e-9/ceil(47.9995e-3)):0))/1)/((((480e-9/ceil(47.9995e-3))*ceil(47.9995e-3))*(480e-9/ceil(47.9995e-3)))*ceil(47.9995e-3))' NRS='480e-9/ceil(47.9995e-3)<119.5e-9?(((14.4e-15+(480e-9/ceil(47.9995e-3))*50e-9)+floor((ceil(47.9995e-3)-1)/2.0)*(14.4e-15+(480e-9/ceil(47.9995e-3))*100e-9))+(ceil(47.9995e-3)/2-floor(ceil(47.9995e-3)/2)==0?14.4e-15+(480e-9/ceil(47.9995e-3))*50e-9:0))/1:(((140e-9*(480e-9/ceil(47.9995e-3))+floor((ceil(47.9995e-3)-1)/2.0)*(110e-9*(480e-9/ceil(47.9995e-3))))+(ceil(47.9995e-3)/2-floor(ceil(47.9995e-3)/2)==0?140e-9*(480e-9/ceil(47.9995e-3)):0))/1)/((((480e-9/ceil(47.9995e-3))*ceil(47.9995e-3))*(480e-9/ceil(47.9995e-3)))*ceil(47.9995e-3))' M=1
.ends level_shifter_1_1_to_1_8
** End of subcircuit definition.

** Library name: ece_482_pdn_v2
** Cell name: unitcell_decap
** View name: schematic
.subckt unitcell_decap vddio vss
m0 net1 net2 vss vss g45n2svt L=150e-9 W=18e-6 AD=1.8e-12 AS=2.1e-12 PD=19.2e-6 PS=25.4e-6 NRD=5.55556e-3 NRS=6.48148e-3 M=1
m1 net2 net1 vddio vddio g45p2svt L=150e-9 W=18e-6 AD=1.8e-12 AS=2.1e-12 PD=19.2e-6 PS=25.4e-6 NRD=5.55556e-3 NRS=6.48148e-3 M=1
.ends unitcell_decap
** End of subcircuit definition.

** Library name: ece_482_pdn_v2
** Cell name: decap3x3x2
** View name: schematic
.subckt decap3x3x2 vddio vss
xi1<0> vddio vss unitcell_decap
xi1<1> vddio vss unitcell_decap
xi1<2> vddio vss unitcell_decap
xi1<3> vddio vss unitcell_decap
xi1<4> vddio vss unitcell_decap
xi1<5> vddio vss unitcell_decap
xi1<6> vddio vss unitcell_decap
xi1<7> vddio vss unitcell_decap
xi1<8> vddio vss unitcell_decap
xi1<9> vddio vss unitcell_decap
xi1<10> vddio vss unitcell_decap
xi1<11> vddio vss unitcell_decap
xi1<12> vddio vss unitcell_decap
xi1<13> vddio vss unitcell_decap
xi1<14> vddio vss unitcell_decap
xi1<15> vddio vss unitcell_decap
xi1<16> vddio vss unitcell_decap
xi1<17> vddio vss unitcell_decap
xi1<18> vddio vss unitcell_decap
xi1<19> vddio vss unitcell_decap
xi1<20> vddio vss unitcell_decap
xi1<21> vddio vss unitcell_decap
xi1<22> vddio vss unitcell_decap
xi1<23> vddio vss unitcell_decap
xi1<24> vddio vss unitcell_decap
xi1<25> vddio vss unitcell_decap
xi1<26> vddio vss unitcell_decap
xi1<27> vddio vss unitcell_decap
xi1<28> vddio vss unitcell_decap
xi1<29> vddio vss unitcell_decap
xi1<30> vddio vss unitcell_decap
xi1<31> vddio vss unitcell_decap
xi1<32> vddio vss unitcell_decap
xi1<33> vddio vss unitcell_decap
xi1<34> vddio vss unitcell_decap
xi1<35> vddio vss unitcell_decap
xi1<36> vddio vss unitcell_decap
xi1<37> vddio vss unitcell_decap
xi1<38> vddio vss unitcell_decap
xi1<39> vddio vss unitcell_decap
.ends decap3x3x2
** End of subcircuit definition.

** Library name: test2
** Cell name: half_adder
** View name: schematic
.subckt half_adder a b c_out s vdd vss
mnm5 vss s c_out vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mnm3 a_xor_b_bar s vss vss g45n1svt L=45e-9 W=480e-9 AD=38.4e-15 AS=52.8e-15 PD=1.12e-6 PS=1.6e-6 NRD=166.667e-3 NRS=229.167e-3 M=1
mnm4 b a_xor_b_bar c_out vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mnm2 s net8 b vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mnm0 s b net8 vss g45n1svt L=45e-9 W=240e-9 AD=19.2e-15 AS=33.6e-15 PD=560e-9 PS=1.04e-6 NRD=333.333e-3 NRS=583.333e-3 M=1
mnm1 net8 a vss vss g45n1svt L=45e-9 W=480e-9 AD=38.4e-15 AS=52.8e-15 PD=1.12e-6 PS=1.6e-6 NRD=166.667e-3 NRS=229.167e-3 M=1
mpm7 b s c_out vdd g45p1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=583.333e-3 NRS=583.333e-3 M=1
mpm5 s a b vdd g45p1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=583.333e-3 NRS=583.333e-3 M=1
mpm8 vss a_xor_b_bar c_out vdd g45p1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=583.333e-3 NRS=583.333e-3 M=1
mpm6 a_xor_b_bar s vdd vdd g45p1svt L=45e-9 W=960e-9 AD=76.8e-15 AS=105.6e-15 PD=1.6e-6 PS=2.32e-6 NRD=83.3333e-3 NRS=114.583e-3 M=1
mpm0 s b a vdd g45p1svt L=45e-9 W=480e-9 AD=38.4e-15 AS=67.2e-15 PD=800e-9 PS=1.52e-6 NRD=166.667e-3 NRS=291.667e-3 M=1
mpm4 net8 a vdd vdd g45p1svt L=45e-9 W=960e-9 AD=76.8e-15 AS=105.6e-15 PD=1.6e-6 PS=2.32e-6 NRD=83.3333e-3 NRS=114.583e-3 M=1
.ends half_adder
** End of subcircuit definition.

** Library name: test2
** Cell name: full_adder
** View name: schematic
.subckt full_adder a b c c_out s vdd vss
mnm6 c a_xor_b_bar s vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mnm4 b a_xor_b_bar c_out vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mnm3 a_xor_b_bar a_xor_b vss vss g45n1svt L=45e-9 W=480e-9 AD=38.4e-15 AS=52.8e-15 PD=1.12e-6 PS=1.6e-6 NRD=166.667e-3 NRS=229.167e-3 M=1
mnm2 net1 c vss vss g45n1svt L=45e-9 W=480e-9 AD=38.4e-15 AS=52.8e-15 PD=1.12e-6 PS=1.6e-6 NRD=166.667e-3 NRS=229.167e-3 M=1
mnm0 a_xor_b b net4 vss g45n1svt L=45e-9 W=240e-9 AD=19.2e-15 AS=33.6e-15 PD=560e-9 PS=1.04e-6 NRD=333.333e-3 NRS=583.333e-3 M=1
mnm1 net4 a vss vss g45n1svt L=45e-9 W=480e-9 AD=38.4e-15 AS=52.8e-15 PD=1.12e-6 PS=1.6e-6 NRD=166.667e-3 NRS=229.167e-3 M=1
mnm8 a_xor_b net4 b vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mnm5 c a_xor_b c_out vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mnm7 net1 a_xor_b s vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
mpm8 a_xor_b a b vdd g45p1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=583.333e-3 NRS=583.333e-3 M=1
mpm7 net1 a_xor_b_bar s vdd g45p1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=583.333e-3 NRS=583.333e-3 M=1
mpm4 b a_xor_b c_out vdd g45p1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=583.333e-3 NRS=583.333e-3 M=1
mpm1 net4 a vdd vdd g45p1svt L=45e-9 W=960e-9 AD=76.8e-15 AS=105.6e-15 PD=1.6e-6 PS=2.32e-6 NRD=83.3333e-3 NRS=114.583e-3 M=1
mpm0 a_xor_b b a vdd g45p1svt L=45e-9 W=480e-9 AD=38.4e-15 AS=67.2e-15 PD=800e-9 PS=1.52e-6 NRD=166.667e-3 NRS=291.667e-3 M=1
mpm2 net1 c vdd vdd g45p1svt L=45e-9 W=960e-9 AD=76.8e-15 AS=105.6e-15 PD=1.6e-6 PS=2.32e-6 NRD=83.3333e-3 NRS=114.583e-3 M=1
mpm3 a_xor_b_bar a_xor_b vdd vdd g45p1svt L=45e-9 W=960e-9 AD=76.8e-15 AS=105.6e-15 PD=1.6e-6 PS=2.32e-6 NRD=83.3333e-3 NRS=114.583e-3 M=1
mpm5 c a_xor_b_bar c_out vdd g45p1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=583.333e-3 NRS=583.333e-3 M=1
mpm6 c a_xor_b s vdd g45p1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=583.333e-3 NRS=583.333e-3 M=1
.ends full_adder
** End of subcircuit definition.

** Library name: test2
** Cell name: inverter_minsize
** View name: schematic
.subckt inverter_minsize in out vdd vss
mpm0 out in vdd vdd g45p1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=583.333e-3 NRS=583.333e-3 M=1
mnm0 out in vss vss g45n1svt L=45e-9 W=120e-9 AD=16.8e-15 AS=16.8e-15 PD=520e-9 PS=520e-9 NRD=1.16667 NRS=1.16667 M=1
.ends inverter_minsize
** End of subcircuit definition.

** Library name: test2
** Cell name: and_minsize
** View name: schematic
.subckt and_minsize a b out vdd vss
mpm1 net1 b vdd vdd g45p1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=583.333e-3 NRS=583.333e-3 M=1
mpm0 net1 a vdd vdd g45p1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=583.333e-3 NRS=583.333e-3 M=1
mnm1 net10 b vss vss g45n1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=583.333e-3 NRS=583.333e-3 M=1
mnm0 net1 a net10 vss g45n1svt L=45e-9 W=240e-9 AD=33.6e-15 AS=33.6e-15 PD=760e-9 PS=760e-9 NRD=583.333e-3 NRS=583.333e-3 M=1
xi0 net1 out vdd vss inverter_minsize
.ends and_minsize
** End of subcircuit definition.

** Library name: test2
** Cell name: level_shifter_1_8_to_1_1
** View name: schematic
.subckt level_shifter_1_8_to_1_1 aio aio_bar a_core a_core_bar vdd vss
m1 a_core aio_bar vss vss g45n2svt L=150e-9 W=640e-9 AD=96e-15 AS=96e-15 PD=1.58e-6 PS=1.58e-6 NRD=234.375e-3 NRS=234.375e-3 M=1
m0 a_core_bar aio vss vss g45n2svt L=150e-9 W=640e-9 AD=96e-15 AS=96e-15 PD=1.58e-6 PS=1.58e-6 NRD=234.375e-3 NRS=234.375e-3 M=1
mpm1 a_core a_core_bar vdd vdd g45p1svt L=45e-9 W=480e-9 AD=67.2e-15 AS=67.2e-15 PD=1.24e-6 PS=1.24e-6 NRD=291.667e-3 NRS=291.667e-3 M=1
mpm0 a_core_bar a_core vdd vdd g45p1svt L=45e-9 W=480e-9 AD=67.2e-15 AS=67.2e-15 PD=1.24e-6 PS=1.24e-6 NRD=291.667e-3 NRS=291.667e-3 M=1
.ends level_shifter_1_8_to_1_1
** End of subcircuit definition.

** Library name: test2
** Cell name: inverter_1_8_v
** View name: schematic
.subckt inverter_1_8_v in out vddio vssio
m0 out in vssio vssio g45n2svt L=150e-9 W=320e-9 AD=48e-15 AS=48e-15 PD=940e-9 PS=940e-9 NRD=468.75e-3 NRS=468.75e-3 M=1
m1 out in vddio vddio g45p2svt L=150e-9 W=640e-9 AD=96e-15 AS=96e-15 PD=1.58e-6 PS=1.58e-6 NRD=234.375e-3 NRS=234.375e-3 M=1
.ends inverter_1_8_v
** End of subcircuit definition.

** Library name: test2
** Cell name: C2MOS_register
** View name: schematic
.subckt C2MOS_register clk clk_bar d q rst vdd vss
mpm3 net17 x vdd vdd g45p1svt L=45e-9 W=240e-9 AD='240e-9/ceil(23.9995e-3)<119.5e-9?(floor(ceil(23.9995e-3)/2.0)*(14.4e-15+(240e-9/ceil(23.9995e-3))*100e-9)+(ceil(23.9995e-3)/2-floor(ceil(23.9995e-3)/2)!=0?14.4e-15+(240e-9/ceil(23.9995e-3))*50e-9:0))/1:(floor(ceil(23.9995e-3)/2.0)*(110e-9*(240e-9/ceil(23.9995e-3)))+(ceil(23.9995e-3)/2-floor(ceil(23.9995e-3)/2)!=0?140e-9*(240e-9/ceil(23.9995e-3)):0))/1' AS='240e-9/ceil(23.9995e-3)<119.5e-9?(((14.4e-15+(240e-9/ceil(23.9995e-3))*50e-9)+floor((ceil(23.9995e-3)-1)/2.0)*(14.4e-15+(240e-9/ceil(23.9995e-3))*100e-9))+(ceil(23.9995e-3)/2-floor(ceil(23.9995e-3)/2)==0?14.4e-15+(240e-9/ceil(23.9995e-3))*50e-9:0))/1:((140e-9*(240e-9/ceil(23.9995e-3))+floor((ceil(23.9995e-3)-1)/2.0)*(110e-9*(240e-9/ceil(23.9995e-3))))+(ceil(23.9995e-3)/2-floor(ceil(23.9995e-3)/2)==0?140e-9*(240e-9/ceil(23.9995e-3)):0))/1'
+PD='240e-9/ceil(23.9995e-3)<119.5e-9?(floor(ceil(23.9995e-3)/2.0)*680e-9+(ceil(23.9995e-3)/2-floor(ceil(23.9995e-3)/2)!=0?580e-9:0))/1:(floor(ceil(23.9995e-3)/2.0)*(220e-9+2*(240e-9/ceil(23.9995e-3)))+(ceil(23.9995e-3)/2-floor(ceil(23.9995e-3)/2)!=0?280e-9+2*(240e-9/ceil(23.9995e-3)):0))/1' PS='240e-9/ceil(23.9995e-3)<119.5e-9?((580e-9+floor((ceil(23.9995e-3)-1)/2.0)*680e-9)+(ceil(23.9995e-3)/2-floor(ceil(23.9995e-3)/2)==0?580e-9:0))/1:(((280e-9+2*(240e-9/ceil(23.9995e-3)))+floor((ceil(23.9995e-3)-1)/2.0)*(220e-9+2*(240e-9/ceil(23.9995e-3))))+(ceil(23.9995e-3)/2-floor(ceil(23.9995e-3)/2)==0?280e-9+2*(240e-9/ceil(23.9995e-3)):0))/1'
+NRD='240e-9/ceil(23.9995e-3)<119.5e-9?(floor(ceil(23.9995e-3)/2.0)*(14.4e-15+(240e-9/ceil(23.9995e-3))*100e-9)+(ceil(23.9995e-3)/2-floor(ceil(23.9995e-3)/2)!=0?14.4e-15+(240e-9/ceil(23.9995e-3))*50e-9:0))/1:((floor(ceil(23.9995e-3)/2.0)*(110e-9*(240e-9/ceil(23.9995e-3)))+(ceil(23.9995e-3)/2-floor(ceil(23.9995e-3)/2)!=0?140e-9*(240e-9/ceil(23.9995e-3)):0))/1)/((((240e-9/ceil(23.9995e-3))*ceil(23.9995e-3))*(240e-9/ceil(23.9995e-3)))*ceil(23.9995e-3))' NRS='240e-9/ceil(23.9995e-3)<119.5e-9?(((14.4e-15+(240e-9/ceil(23.9995e-3))*50e-9)+floor((ceil(23.9995e-3)-1)/2.0)*(14.4e-15+(240e-9/ceil(23.9995e-3))*100e-9))+(ceil(23.9995e-3)/2-floor(ceil(23.9995e-3)/2)==0?14.4e-15+(240e-9/ceil(23.9995e-3))*50e-9:0))/1:(((140e-9*(240e-9/ceil(23.9995e-3))+floor((ceil(23.9995e-3)-1)/2.0)*(110e-9*(240e-9/ceil(23.9995e-3))))+(ceil(23.9995e-3)/2-floor(ceil(23.9995e-3)/2)==0?140e-9*(240e-9/ceil(23.9995e-3)):0))/1)/((((240e-9/ceil(23.9995e-3))*ceil(23.9995e-3))*(240e-9/ceil(23.9995e-3)))*ceil(23.9995e-3))' M=1
mpm2 q clk_bar net17 vdd g45p1svt L=45e-9 W=240e-9 AD='240e-9/ceil(23.9995e-3)<119.5e-9?(floor(ceil(23.9995e-3)/2.0)*(14.4e-15+(240e-9/ceil(23.9995e-3))*100e-9)+(ceil(23.9995e-3)/2-floor(ceil(23.9995e-3)/2)!=0?14.4e-15+(240e-9/ceil(23.9995e-3))*50e-9:0))/1:(floor(ceil(23.9995e-3)/2.0)*(110e-9*(240e-9/ceil(23.9995e-3)))+(ceil(23.9995e-3)/2-floor(ceil(23.9995e-3)/2)!=0?140e-9*(240e-9/ceil(23.9995e-3)):0))/1' AS='240e-9/ceil(23.9995e-3)<119.5e-9?(((14.4e-15+(240e-9/ceil(23.9995e-3))*50e-9)+floor((ceil(23.9995e-3)-1)/2.0)*(14.4e-15+(240e-9/ceil(23.9995e-3))*100e-9))+(ceil(23.9995e-3)/2-floor(ceil(23.9995e-3)/2)==0?14.4e-15+(240e-9/ceil(23.9995e-3))*50e-9:0))/1:((140e-9*(240e-9/ceil(23.9995e-3))+floor((ceil(23.9995e-3)-1)/2.0)*(110e-9*(240e-9/ceil(23.9995e-3))))+(ceil(23.9995e-3)/2-floor(ceil(23.9995e-3)/2)==0?140e-9*(240e-9/ceil(23.9995e-3)):0))/1'
+PD='240e-9/ceil(23.9995e-3)<119.5e-9?(floor(ceil(23.9995e-3)/2.0)*680e-9+(ceil(23.9995e-3)/2-floor(ceil(23.9995e-3)/2)!=0?580e-9:0))/1:(floor(ceil(23.9995e-3)/2.0)*(220e-9+2*(240e-9/ceil(23.9995e-3)))+(ceil(23.9995e-3)/2-floor(ceil(23.9995e-3)/2)!=0?280e-9+2*(240e-9/ceil(23.9995e-3)):0))/1' PS='240e-9/ceil(23.9995e-3)<119.5e-9?((580e-9+floor((ceil(23.9995e-3)-1)/2.0)*680e-9)+(ceil(23.9995e-3)/2-floor(ceil(23.9995e-3)/2)==0?580e-9:0))/1:(((280e-9+2*(240e-9/ceil(23.9995e-3)))+floor((ceil(23.9995e-3)-1)/2.0)*(220e-9+2*(240e-9/ceil(23.9995e-3))))+(ceil(23.9995e-3)/2-floor(ceil(23.9995e-3)/2)==0?280e-9+2*(240e-9/ceil(23.9995e-3)):0))/1'
+NRD='240e-9/ceil(23.9995e-3)<119.5e-9?(floor(ceil(23.9995e-3)/2.0)*(14.4e-15+(240e-9/ceil(23.9995e-3))*100e-9)+(ceil(23.9995e-3)/2-floor(ceil(23.9995e-3)/2)!=0?14.4e-15+(240e-9/ceil(23.9995e-3))*50e-9:0))/1:((floor(ceil(23.9995e-3)/2.0)*(110e-9*(240e-9/ceil(23.9995e-3)))+(ceil(23.9995e-3)/2-floor(ceil(23.9995e-3)/2)!=0?140e-9*(240e-9/ceil(23.9995e-3)):0))/1)/((((240e-9/ceil(23.9995e-3))*ceil(23.9995e-3))*(240e-9/ceil(23.9995e-3)))*ceil(23.9995e-3))' NRS='240e-9/ceil(23.9995e-3)<119.5e-9?(((14.4e-15+(240e-9/ceil(23.9995e-3))*50e-9)+floor((ceil(23.9995e-3)-1)/2.0)*(14.4e-15+(240e-9/ceil(23.9995e-3))*100e-9))+(ceil(23.9995e-3)/2-floor(ceil(23.9995e-3)/2)==0?14.4e-15+(240e-9/ceil(23.9995e-3))*50e-9:0))/1:(((140e-9*(240e-9/ceil(23.9995e-3))+floor((ceil(23.9995e-3)-1)/2.0)*(110e-9*(240e-9/ceil(23.9995e-3))))+(ceil(23.9995e-3)/2-floor(ceil(23.9995e-3)/2)==0?140e-9*(240e-9/ceil(23.9995e-3)):0))/1)/((((240e-9/ceil(23.9995e-3))*ceil(23.9995e-3))*(240e-9/ceil(23.9995e-3)))*ceil(23.9995e-3))' M=1
mpm1 x clk net4 vdd g45p1svt L=45e-9 W=240e-9 AD='240e-9/ceil(23.9995e-3)<119.5e-9?(floor(ceil(23.9995e-3)/2.0)*(14.4e-15+(240e-9/ceil(23.9995e-3))*100e-9)+(ceil(23.9995e-3)/2-floor(ceil(23.9995e-3)/2)!=0?14.4e-15+(240e-9/ceil(23.9995e-3))*50e-9:0))/1:(floor(ceil(23.9995e-3)/2.0)*(110e-9*(240e-9/ceil(23.9995e-3)))+(ceil(23.9995e-3)/2-floor(ceil(23.9995e-3)/2)!=0?140e-9*(240e-9/ceil(23.9995e-3)):0))/1' AS='240e-9/ceil(23.9995e-3)<119.5e-9?(((14.4e-15+(240e-9/ceil(23.9995e-3))*50e-9)+floor((ceil(23.9995e-3)-1)/2.0)*(14.4e-15+(240e-9/ceil(23.9995e-3))*100e-9))+(ceil(23.9995e-3)/2-floor(ceil(23.9995e-3)/2)==0?14.4e-15+(240e-9/ceil(23.9995e-3))*50e-9:0))/1:((140e-9*(240e-9/ceil(23.9995e-3))+floor((ceil(23.9995e-3)-1)/2.0)*(110e-9*(240e-9/ceil(23.9995e-3))))+(ceil(23.9995e-3)/2-floor(ceil(23.9995e-3)/2)==0?140e-9*(240e-9/ceil(23.9995e-3)):0))/1'
+PD='240e-9/ceil(23.9995e-3)<119.5e-9?(floor(ceil(23.9995e-3)/2.0)*680e-9+(ceil(23.9995e-3)/2-floor(ceil(23.9995e-3)/2)!=0?580e-9:0))/1:(floor(ceil(23.9995e-3)/2.0)*(220e-9+2*(240e-9/ceil(23.9995e-3)))+(ceil(23.9995e-3)/2-floor(ceil(23.9995e-3)/2)!=0?280e-9+2*(240e-9/ceil(23.9995e-3)):0))/1' PS='240e-9/ceil(23.9995e-3)<119.5e-9?((580e-9+floor((ceil(23.9995e-3)-1)/2.0)*680e-9)+(ceil(23.9995e-3)/2-floor(ceil(23.9995e-3)/2)==0?580e-9:0))/1:(((280e-9+2*(240e-9/ceil(23.9995e-3)))+floor((ceil(23.9995e-3)-1)/2.0)*(220e-9+2*(240e-9/ceil(23.9995e-3))))+(ceil(23.9995e-3)/2-floor(ceil(23.9995e-3)/2)==0?280e-9+2*(240e-9/ceil(23.9995e-3)):0))/1'
+NRD='240e-9/ceil(23.9995e-3)<119.5e-9?(floor(ceil(23.9995e-3)/2.0)*(14.4e-15+(240e-9/ceil(23.9995e-3))*100e-9)+(ceil(23.9995e-3)/2-floor(ceil(23.9995e-3)/2)!=0?14.4e-15+(240e-9/ceil(23.9995e-3))*50e-9:0))/1:((floor(ceil(23.9995e-3)/2.0)*(110e-9*(240e-9/ceil(23.9995e-3)))+(ceil(23.9995e-3)/2-floor(ceil(23.9995e-3)/2)!=0?140e-9*(240e-9/ceil(23.9995e-3)):0))/1)/((((240e-9/ceil(23.9995e-3))*ceil(23.9995e-3))*(240e-9/ceil(23.9995e-3)))*ceil(23.9995e-3))' NRS='240e-9/ceil(23.9995e-3)<119.5e-9?(((14.4e-15+(240e-9/ceil(23.9995e-3))*50e-9)+floor((ceil(23.9995e-3)-1)/2.0)*(14.4e-15+(240e-9/ceil(23.9995e-3))*100e-9))+(ceil(23.9995e-3)/2-floor(ceil(23.9995e-3)/2)==0?14.4e-15+(240e-9/ceil(23.9995e-3))*50e-9:0))/1:(((140e-9*(240e-9/ceil(23.9995e-3))+floor((ceil(23.9995e-3)-1)/2.0)*(110e-9*(240e-9/ceil(23.9995e-3))))+(ceil(23.9995e-3)/2-floor(ceil(23.9995e-3)/2)==0?140e-9*(240e-9/ceil(23.9995e-3)):0))/1)/((((240e-9/ceil(23.9995e-3))*ceil(23.9995e-3))*(240e-9/ceil(23.9995e-3)))*ceil(23.9995e-3))' M=1
mpm0 net4 net5 vdd vdd g45p1svt L=45e-9 W=240e-9 AD='240e-9/ceil(23.9995e-3)<119.5e-9?(floor(ceil(23.9995e-3)/2.0)*(14.4e-15+(240e-9/ceil(23.9995e-3))*100e-9)+(ceil(23.9995e-3)/2-floor(ceil(23.9995e-3)/2)!=0?14.4e-15+(240e-9/ceil(23.9995e-3))*50e-9:0))/1:(floor(ceil(23.9995e-3)/2.0)*(110e-9*(240e-9/ceil(23.9995e-3)))+(ceil(23.9995e-3)/2-floor(ceil(23.9995e-3)/2)!=0?140e-9*(240e-9/ceil(23.9995e-3)):0))/1' AS='240e-9/ceil(23.9995e-3)<119.5e-9?(((14.4e-15+(240e-9/ceil(23.9995e-3))*50e-9)+floor((ceil(23.9995e-3)-1)/2.0)*(14.4e-15+(240e-9/ceil(23.9995e-3))*100e-9))+(ceil(23.9995e-3)/2-floor(ceil(23.9995e-3)/2)==0?14.4e-15+(240e-9/ceil(23.9995e-3))*50e-9:0))/1:((140e-9*(240e-9/ceil(23.9995e-3))+floor((ceil(23.9995e-3)-1)/2.0)*(110e-9*(240e-9/ceil(23.9995e-3))))+(ceil(23.9995e-3)/2-floor(ceil(23.9995e-3)/2)==0?140e-9*(240e-9/ceil(23.9995e-3)):0))/1'
+PD='240e-9/ceil(23.9995e-3)<119.5e-9?(floor(ceil(23.9995e-3)/2.0)*680e-9+(ceil(23.9995e-3)/2-floor(ceil(23.9995e-3)/2)!=0?580e-9:0))/1:(floor(ceil(23.9995e-3)/2.0)*(220e-9+2*(240e-9/ceil(23.9995e-3)))+(ceil(23.9995e-3)/2-floor(ceil(23.9995e-3)/2)!=0?280e-9+2*(240e-9/ceil(23.9995e-3)):0))/1' PS='240e-9/ceil(23.9995e-3)<119.5e-9?((580e-9+floor((ceil(23.9995e-3)-1)/2.0)*680e-9)+(ceil(23.9995e-3)/2-floor(ceil(23.9995e-3)/2)==0?580e-9:0))/1:(((280e-9+2*(240e-9/ceil(23.9995e-3)))+floor((ceil(23.9995e-3)-1)/2.0)*(220e-9+2*(240e-9/ceil(23.9995e-3))))+(ceil(23.9995e-3)/2-floor(ceil(23.9995e-3)/2)==0?280e-9+2*(240e-9/ceil(23.9995e-3)):0))/1'
+NRD='240e-9/ceil(23.9995e-3)<119.5e-9?(floor(ceil(23.9995e-3)/2.0)*(14.4e-15+(240e-9/ceil(23.9995e-3))*100e-9)+(ceil(23.9995e-3)/2-floor(ceil(23.9995e-3)/2)!=0?14.4e-15+(240e-9/ceil(23.9995e-3))*50e-9:0))/1:((floor(ceil(23.9995e-3)/2.0)*(110e-9*(240e-9/ceil(23.9995e-3)))+(ceil(23.9995e-3)/2-floor(ceil(23.9995e-3)/2)!=0?140e-9*(240e-9/ceil(23.9995e-3)):0))/1)/((((240e-9/ceil(23.9995e-3))*ceil(23.9995e-3))*(240e-9/ceil(23.9995e-3)))*ceil(23.9995e-3))' NRS='240e-9/ceil(23.9995e-3)<119.5e-9?(((14.4e-15+(240e-9/ceil(23.9995e-3))*50e-9)+floor((ceil(23.9995e-3)-1)/2.0)*(14.4e-15+(240e-9/ceil(23.9995e-3))*100e-9))+(ceil(23.9995e-3)/2-floor(ceil(23.9995e-3)/2)==0?14.4e-15+(240e-9/ceil(23.9995e-3))*50e-9:0))/1:(((140e-9*(240e-9/ceil(23.9995e-3))+floor((ceil(23.9995e-3)-1)/2.0)*(110e-9*(240e-9/ceil(23.9995e-3))))+(ceil(23.9995e-3)/2-floor(ceil(23.9995e-3)/2)==0?140e-9*(240e-9/ceil(23.9995e-3)):0))/1)/((((240e-9/ceil(23.9995e-3))*ceil(23.9995e-3))*(240e-9/ceil(23.9995e-3)))*ceil(23.9995e-3))' M=1
mnm3 net21 x vss vss g45n1svt L=45e-9 W=120e-9 AD='120e-9/ceil(11.9995e-3)<119.5e-9?(floor(ceil(11.9995e-3)/2.0)*(14.4e-15+(120e-9/ceil(11.9995e-3))*100e-9)+(ceil(11.9995e-3)/2-floor(ceil(11.9995e-3)/2)!=0?14.4e-15+(120e-9/ceil(11.9995e-3))*50e-9:0))/1:(floor(ceil(11.9995e-3)/2.0)*(110e-9*(120e-9/ceil(11.9995e-3)))+(ceil(11.9995e-3)/2-floor(ceil(11.9995e-3)/2)!=0?140e-9*(120e-9/ceil(11.9995e-3)):0))/1' AS='120e-9/ceil(11.9995e-3)<119.5e-9?(((14.4e-15+(120e-9/ceil(11.9995e-3))*50e-9)+floor((ceil(11.9995e-3)-1)/2.0)*(14.4e-15+(120e-9/ceil(11.9995e-3))*100e-9))+(ceil(11.9995e-3)/2-floor(ceil(11.9995e-3)/2)==0?14.4e-15+(120e-9/ceil(11.9995e-3))*50e-9:0))/1:((140e-9*(120e-9/ceil(11.9995e-3))+floor((ceil(11.9995e-3)-1)/2.0)*(110e-9*(120e-9/ceil(11.9995e-3))))+(ceil(11.9995e-3)/2-floor(ceil(11.9995e-3)/2)==0?140e-9*(120e-9/ceil(11.9995e-3)):0))/1'
+PD='120e-9/ceil(11.9995e-3)<119.5e-9?(floor(ceil(11.9995e-3)/2.0)*680e-9+(ceil(11.9995e-3)/2-floor(ceil(11.9995e-3)/2)!=0?580e-9:0))/1:(floor(ceil(11.9995e-3)/2.0)*(220e-9+2*(120e-9/ceil(11.9995e-3)))+(ceil(11.9995e-3)/2-floor(ceil(11.9995e-3)/2)!=0?280e-9+2*(120e-9/ceil(11.9995e-3)):0))/1' PS='120e-9/ceil(11.9995e-3)<119.5e-9?((580e-9+floor((ceil(11.9995e-3)-1)/2.0)*680e-9)+(ceil(11.9995e-3)/2-floor(ceil(11.9995e-3)/2)==0?580e-9:0))/1:(((280e-9+2*(120e-9/ceil(11.9995e-3)))+floor((ceil(11.9995e-3)-1)/2.0)*(220e-9+2*(120e-9/ceil(11.9995e-3))))+(ceil(11.9995e-3)/2-floor(ceil(11.9995e-3)/2)==0?280e-9+2*(120e-9/ceil(11.9995e-3)):0))/1'
+NRD='120e-9/ceil(11.9995e-3)<119.5e-9?(floor(ceil(11.9995e-3)/2.0)*(14.4e-15+(120e-9/ceil(11.9995e-3))*100e-9)+(ceil(11.9995e-3)/2-floor(ceil(11.9995e-3)/2)!=0?14.4e-15+(120e-9/ceil(11.9995e-3))*50e-9:0))/1:((floor(ceil(11.9995e-3)/2.0)*(110e-9*(120e-9/ceil(11.9995e-3)))+(ceil(11.9995e-3)/2-floor(ceil(11.9995e-3)/2)!=0?140e-9*(120e-9/ceil(11.9995e-3)):0))/1)/((((120e-9/ceil(11.9995e-3))*ceil(11.9995e-3))*(120e-9/ceil(11.9995e-3)))*ceil(11.9995e-3))' NRS='120e-9/ceil(11.9995e-3)<119.5e-9?(((14.4e-15+(120e-9/ceil(11.9995e-3))*50e-9)+floor((ceil(11.9995e-3)-1)/2.0)*(14.4e-15+(120e-9/ceil(11.9995e-3))*100e-9))+(ceil(11.9995e-3)/2-floor(ceil(11.9995e-3)/2)==0?14.4e-15+(120e-9/ceil(11.9995e-3))*50e-9:0))/1:(((140e-9*(120e-9/ceil(11.9995e-3))+floor((ceil(11.9995e-3)-1)/2.0)*(110e-9*(120e-9/ceil(11.9995e-3))))+(ceil(11.9995e-3)/2-floor(ceil(11.9995e-3)/2)==0?140e-9*(120e-9/ceil(11.9995e-3)):0))/1)/((((120e-9/ceil(11.9995e-3))*ceil(11.9995e-3))*(120e-9/ceil(11.9995e-3)))*ceil(11.9995e-3))' M=1
mnm2 q clk net21 vss g45n1svt L=45e-9 W=120e-9 AD='120e-9/ceil(11.9995e-3)<119.5e-9?(floor(ceil(11.9995e-3)/2.0)*(14.4e-15+(120e-9/ceil(11.9995e-3))*100e-9)+(ceil(11.9995e-3)/2-floor(ceil(11.9995e-3)/2)!=0?14.4e-15+(120e-9/ceil(11.9995e-3))*50e-9:0))/1:(floor(ceil(11.9995e-3)/2.0)*(110e-9*(120e-9/ceil(11.9995e-3)))+(ceil(11.9995e-3)/2-floor(ceil(11.9995e-3)/2)!=0?140e-9*(120e-9/ceil(11.9995e-3)):0))/1' AS='120e-9/ceil(11.9995e-3)<119.5e-9?(((14.4e-15+(120e-9/ceil(11.9995e-3))*50e-9)+floor((ceil(11.9995e-3)-1)/2.0)*(14.4e-15+(120e-9/ceil(11.9995e-3))*100e-9))+(ceil(11.9995e-3)/2-floor(ceil(11.9995e-3)/2)==0?14.4e-15+(120e-9/ceil(11.9995e-3))*50e-9:0))/1:((140e-9*(120e-9/ceil(11.9995e-3))+floor((ceil(11.9995e-3)-1)/2.0)*(110e-9*(120e-9/ceil(11.9995e-3))))+(ceil(11.9995e-3)/2-floor(ceil(11.9995e-3)/2)==0?140e-9*(120e-9/ceil(11.9995e-3)):0))/1'
+PD='120e-9/ceil(11.9995e-3)<119.5e-9?(floor(ceil(11.9995e-3)/2.0)*680e-9+(ceil(11.9995e-3)/2-floor(ceil(11.9995e-3)/2)!=0?580e-9:0))/1:(floor(ceil(11.9995e-3)/2.0)*(220e-9+2*(120e-9/ceil(11.9995e-3)))+(ceil(11.9995e-3)/2-floor(ceil(11.9995e-3)/2)!=0?280e-9+2*(120e-9/ceil(11.9995e-3)):0))/1' PS='120e-9/ceil(11.9995e-3)<119.5e-9?((580e-9+floor((ceil(11.9995e-3)-1)/2.0)*680e-9)+(ceil(11.9995e-3)/2-floor(ceil(11.9995e-3)/2)==0?580e-9:0))/1:(((280e-9+2*(120e-9/ceil(11.9995e-3)))+floor((ceil(11.9995e-3)-1)/2.0)*(220e-9+2*(120e-9/ceil(11.9995e-3))))+(ceil(11.9995e-3)/2-floor(ceil(11.9995e-3)/2)==0?280e-9+2*(120e-9/ceil(11.9995e-3)):0))/1'
+NRD='120e-9/ceil(11.9995e-3)<119.5e-9?(floor(ceil(11.9995e-3)/2.0)*(14.4e-15+(120e-9/ceil(11.9995e-3))*100e-9)+(ceil(11.9995e-3)/2-floor(ceil(11.9995e-3)/2)!=0?14.4e-15+(120e-9/ceil(11.9995e-3))*50e-9:0))/1:((floor(ceil(11.9995e-3)/2.0)*(110e-9*(120e-9/ceil(11.9995e-3)))+(ceil(11.9995e-3)/2-floor(ceil(11.9995e-3)/2)!=0?140e-9*(120e-9/ceil(11.9995e-3)):0))/1)/((((120e-9/ceil(11.9995e-3))*ceil(11.9995e-3))*(120e-9/ceil(11.9995e-3)))*ceil(11.9995e-3))' NRS='120e-9/ceil(11.9995e-3)<119.5e-9?(((14.4e-15+(120e-9/ceil(11.9995e-3))*50e-9)+floor((ceil(11.9995e-3)-1)/2.0)*(14.4e-15+(120e-9/ceil(11.9995e-3))*100e-9))+(ceil(11.9995e-3)/2-floor(ceil(11.9995e-3)/2)==0?14.4e-15+(120e-9/ceil(11.9995e-3))*50e-9:0))/1:(((140e-9*(120e-9/ceil(11.9995e-3))+floor((ceil(11.9995e-3)-1)/2.0)*(110e-9*(120e-9/ceil(11.9995e-3))))+(ceil(11.9995e-3)/2-floor(ceil(11.9995e-3)/2)==0?140e-9*(120e-9/ceil(11.9995e-3)):0))/1)/((((120e-9/ceil(11.9995e-3))*ceil(11.9995e-3))*(120e-9/ceil(11.9995e-3)))*ceil(11.9995e-3))' M=1
mnm1 net9 net5 vss vss g45n1svt L=45e-9 W=120e-9 AD='120e-9/ceil(11.9995e-3)<119.5e-9?(floor(ceil(11.9995e-3)/2.0)*(14.4e-15+(120e-9/ceil(11.9995e-3))*100e-9)+(ceil(11.9995e-3)/2-floor(ceil(11.9995e-3)/2)!=0?14.4e-15+(120e-9/ceil(11.9995e-3))*50e-9:0))/1:(floor(ceil(11.9995e-3)/2.0)*(110e-9*(120e-9/ceil(11.9995e-3)))+(ceil(11.9995e-3)/2-floor(ceil(11.9995e-3)/2)!=0?140e-9*(120e-9/ceil(11.9995e-3)):0))/1' AS='120e-9/ceil(11.9995e-3)<119.5e-9?(((14.4e-15+(120e-9/ceil(11.9995e-3))*50e-9)+floor((ceil(11.9995e-3)-1)/2.0)*(14.4e-15+(120e-9/ceil(11.9995e-3))*100e-9))+(ceil(11.9995e-3)/2-floor(ceil(11.9995e-3)/2)==0?14.4e-15+(120e-9/ceil(11.9995e-3))*50e-9:0))/1:((140e-9*(120e-9/ceil(11.9995e-3))+floor((ceil(11.9995e-3)-1)/2.0)*(110e-9*(120e-9/ceil(11.9995e-3))))+(ceil(11.9995e-3)/2-floor(ceil(11.9995e-3)/2)==0?140e-9*(120e-9/ceil(11.9995e-3)):0))/1'
+PD='120e-9/ceil(11.9995e-3)<119.5e-9?(floor(ceil(11.9995e-3)/2.0)*680e-9+(ceil(11.9995e-3)/2-floor(ceil(11.9995e-3)/2)!=0?580e-9:0))/1:(floor(ceil(11.9995e-3)/2.0)*(220e-9+2*(120e-9/ceil(11.9995e-3)))+(ceil(11.9995e-3)/2-floor(ceil(11.9995e-3)/2)!=0?280e-9+2*(120e-9/ceil(11.9995e-3)):0))/1' PS='120e-9/ceil(11.9995e-3)<119.5e-9?((580e-9+floor((ceil(11.9995e-3)-1)/2.0)*680e-9)+(ceil(11.9995e-3)/2-floor(ceil(11.9995e-3)/2)==0?580e-9:0))/1:(((280e-9+2*(120e-9/ceil(11.9995e-3)))+floor((ceil(11.9995e-3)-1)/2.0)*(220e-9+2*(120e-9/ceil(11.9995e-3))))+(ceil(11.9995e-3)/2-floor(ceil(11.9995e-3)/2)==0?280e-9+2*(120e-9/ceil(11.9995e-3)):0))/1'
+NRD='120e-9/ceil(11.9995e-3)<119.5e-9?(floor(ceil(11.9995e-3)/2.0)*(14.4e-15+(120e-9/ceil(11.9995e-3))*100e-9)+(ceil(11.9995e-3)/2-floor(ceil(11.9995e-3)/2)!=0?14.4e-15+(120e-9/ceil(11.9995e-3))*50e-9:0))/1:((floor(ceil(11.9995e-3)/2.0)*(110e-9*(120e-9/ceil(11.9995e-3)))+(ceil(11.9995e-3)/2-floor(ceil(11.9995e-3)/2)!=0?140e-9*(120e-9/ceil(11.9995e-3)):0))/1)/((((120e-9/ceil(11.9995e-3))*ceil(11.9995e-3))*(120e-9/ceil(11.9995e-3)))*ceil(11.9995e-3))' NRS='120e-9/ceil(11.9995e-3)<119.5e-9?(((14.4e-15+(120e-9/ceil(11.9995e-3))*50e-9)+floor((ceil(11.9995e-3)-1)/2.0)*(14.4e-15+(120e-9/ceil(11.9995e-3))*100e-9))+(ceil(11.9995e-3)/2-floor(ceil(11.9995e-3)/2)==0?14.4e-15+(120e-9/ceil(11.9995e-3))*50e-9:0))/1:(((140e-9*(120e-9/ceil(11.9995e-3))+floor((ceil(11.9995e-3)-1)/2.0)*(110e-9*(120e-9/ceil(11.9995e-3))))+(ceil(11.9995e-3)/2-floor(ceil(11.9995e-3)/2)==0?140e-9*(120e-9/ceil(11.9995e-3)):0))/1)/((((120e-9/ceil(11.9995e-3))*ceil(11.9995e-3))*(120e-9/ceil(11.9995e-3)))*ceil(11.9995e-3))' M=1
mnm0 x clk_bar net9 vss g45n1svt L=45e-9 W=120e-9 AD='120e-9/ceil(11.9995e-3)<119.5e-9?(floor(ceil(11.9995e-3)/2.0)*(14.4e-15+(120e-9/ceil(11.9995e-3))*100e-9)+(ceil(11.9995e-3)/2-floor(ceil(11.9995e-3)/2)!=0?14.4e-15+(120e-9/ceil(11.9995e-3))*50e-9:0))/1:(floor(ceil(11.9995e-3)/2.0)*(110e-9*(120e-9/ceil(11.9995e-3)))+(ceil(11.9995e-3)/2-floor(ceil(11.9995e-3)/2)!=0?140e-9*(120e-9/ceil(11.9995e-3)):0))/1' AS='120e-9/ceil(11.9995e-3)<119.5e-9?(((14.4e-15+(120e-9/ceil(11.9995e-3))*50e-9)+floor((ceil(11.9995e-3)-1)/2.0)*(14.4e-15+(120e-9/ceil(11.9995e-3))*100e-9))+(ceil(11.9995e-3)/2-floor(ceil(11.9995e-3)/2)==0?14.4e-15+(120e-9/ceil(11.9995e-3))*50e-9:0))/1:((140e-9*(120e-9/ceil(11.9995e-3))+floor((ceil(11.9995e-3)-1)/2.0)*(110e-9*(120e-9/ceil(11.9995e-3))))+(ceil(11.9995e-3)/2-floor(ceil(11.9995e-3)/2)==0?140e-9*(120e-9/ceil(11.9995e-3)):0))/1'
+PD='120e-9/ceil(11.9995e-3)<119.5e-9?(floor(ceil(11.9995e-3)/2.0)*680e-9+(ceil(11.9995e-3)/2-floor(ceil(11.9995e-3)/2)!=0?580e-9:0))/1:(floor(ceil(11.9995e-3)/2.0)*(220e-9+2*(120e-9/ceil(11.9995e-3)))+(ceil(11.9995e-3)/2-floor(ceil(11.9995e-3)/2)!=0?280e-9+2*(120e-9/ceil(11.9995e-3)):0))/1' PS='120e-9/ceil(11.9995e-3)<119.5e-9?((580e-9+floor((ceil(11.9995e-3)-1)/2.0)*680e-9)+(ceil(11.9995e-3)/2-floor(ceil(11.9995e-3)/2)==0?580e-9:0))/1:(((280e-9+2*(120e-9/ceil(11.9995e-3)))+floor((ceil(11.9995e-3)-1)/2.0)*(220e-9+2*(120e-9/ceil(11.9995e-3))))+(ceil(11.9995e-3)/2-floor(ceil(11.9995e-3)/2)==0?280e-9+2*(120e-9/ceil(11.9995e-3)):0))/1'
+NRD='120e-9/ceil(11.9995e-3)<119.5e-9?(floor(ceil(11.9995e-3)/2.0)*(14.4e-15+(120e-9/ceil(11.9995e-3))*100e-9)+(ceil(11.9995e-3)/2-floor(ceil(11.9995e-3)/2)!=0?14.4e-15+(120e-9/ceil(11.9995e-3))*50e-9:0))/1:((floor(ceil(11.9995e-3)/2.0)*(110e-9*(120e-9/ceil(11.9995e-3)))+(ceil(11.9995e-3)/2-floor(ceil(11.9995e-3)/2)!=0?140e-9*(120e-9/ceil(11.9995e-3)):0))/1)/((((120e-9/ceil(11.9995e-3))*ceil(11.9995e-3))*(120e-9/ceil(11.9995e-3)))*ceil(11.9995e-3))' NRS='120e-9/ceil(11.9995e-3)<119.5e-9?(((14.4e-15+(120e-9/ceil(11.9995e-3))*50e-9)+floor((ceil(11.9995e-3)-1)/2.0)*(14.4e-15+(120e-9/ceil(11.9995e-3))*100e-9))+(ceil(11.9995e-3)/2-floor(ceil(11.9995e-3)/2)==0?14.4e-15+(120e-9/ceil(11.9995e-3))*50e-9:0))/1:(((140e-9*(120e-9/ceil(11.9995e-3))+floor((ceil(11.9995e-3)-1)/2.0)*(110e-9*(120e-9/ceil(11.9995e-3))))+(ceil(11.9995e-3)/2-floor(ceil(11.9995e-3)/2)==0?140e-9*(120e-9/ceil(11.9995e-3)):0))/1)/((((120e-9/ceil(11.9995e-3))*ceil(11.9995e-3))*(120e-9/ceil(11.9995e-3)))*ceil(11.9995e-3))' M=1
xi0 d net8 net5 vdd vss and_minsize
xi1 rst net8 vdd vss inverter_minsize
.ends C2MOS_register
** End of subcircuit definition.

** Library name: test2
** Cell name: superbuffer_4
** View name: schematic
.subckt superbuffer_4 vddio vss sbuf_in sbuf_out
m7 net17 net7 vddio vddio g45p2svt L=150e-9 W=40.96e-6 AD=4.50725e-12 AS=4.50725e-12 PD=50.27e-6 PS=50.27e-6 NRD=2.68456e-3 NRS=2.68456e-3 M=1
m4 sbuf_out net17 vddio vddio g45p2svt L=150e-9 W=163.84e-6 AD=16.87e-12 AS=16.87e-12 PD=177.02e-6 PS=177.02e-6 NRD=628.15e-6 NRS=628.15e-6 M=1
m1 net7 net3 vddio vddio g45p2svt L=150e-9 W=10.24e-6 AD=1.024e-12 AS=1.28e-12 PD=11.04e-6 PS=16.36e-6 NRD=9.76562e-3 NRS=12.207e-3 M=1
m0 net3 sbuf_in vddio vddio g45p2svt L=150e-9 W=2.56e-6 AD=384e-15 AS=384e-15 PD=5.42e-6 PS=5.42e-6 NRD=58.5937e-3 NRS=58.5937e-3 M=1
m6 sbuf_out net17 vss vss g45n2svt L=150e-9 W=81.92e-6 AD=8.192e-12 AS=8.704e-12 PD=85.12e-6 PS=95.56e-6 NRD=1.2207e-3 NRS=1.297e-3 M=1
m5 net17 net7 vss vss g45n2svt L=150e-9 W=20.48e-6 AD=2.048e-12 AS=2.56e-12 PD=21.28e-6 PS=31.72e-6 NRD=4.88281e-3 NRS=6.10352e-3 M=1
m3 net7 net3 vss vss g45n2svt L=150e-9 W=5.12e-6 AD=512e-15 AS=640e-15 PD=5.92e-6 PS=8.68e-6 NRD=19.5312e-3 NRS=24.4141e-3 M=1
m2 net3 sbuf_in vss vss g45n2svt L=150e-9 W=1.28e-6 AD=192e-15 AS=192e-15 PD=2.86e-6 PS=2.86e-6 NRD=117.187e-3 NRS=117.187e-3 M=1
.ends superbuffer_4
** End of subcircuit definition.

** Library name: test2
** Cell name: multiplier
** View name: schematic
xi117 p7_f p7_bar p7_1_1 net59 vddio1 vss1 level_shifter_1_1_to_1_8
xi116 p6_f p6_bar p6_1_1 net53 vddio1 vss1 level_shifter_1_1_to_1_8
xi115 p5_f p5_bar p5_1_1 net47 vddio1 vss1 level_shifter_1_1_to_1_8
xi114 p4_f p4_bar p4_1_1 net38 vddio1 vss1 level_shifter_1_1_to_1_8
xi113 p3_f p3_bar p3_1_1 net30 vddio1 vss1 level_shifter_1_1_to_1_8
xi112 p2_f p2_bar p2_1_1 net24 vddio1 vss1 level_shifter_1_1_to_1_8
xi111 p1_f p1_bar p1_1_1 net16 vddio1 vss1 level_shifter_1_1_to_1_8
xi110 p0_f p0_bar p0_1_1 net7 vddio1 vss1 level_shifter_1_1_to_1_8
xi126 vddio1 vss1 decap3x3x2
xi133 vddio1 vss1 decap3x3x2
xi134 vddio1 vss1 decap3x3x2
xi131 vddio1 vss1 decap3x3x2
xi132 vddio1 vss1 decap3x3x2
xi130 vddio1 vss1 decap3x3x2
xi129 vddio1 vss1 decap3x3x2
xi128 vddio1 vss1 decap3x3x2
xi127 vddio1 vss1 decap3x3x2
xi29 s_1_1_reg net6 c_2_0 p_3 vdd1 vss1 half_adder
xi20 s_0_1_reg net5 c_1_0 p_2 vdd1 vss1 half_adder
xi15 c_0_2 net41 c_0_3 s_0_3 vdd1 vss1 half_adder
xi137 net10 net8 c_0_0 p_1 vdd1 vss1 half_adder
xi32 c_1_3_reg net11 c_2_2 p_7 p_6 vdd1 vss1 full_adder
xi31 s_1_3_reg net1 c_2_1 c_2_2 p_5 vdd1 vss1 full_adder
xi30 s_1_2_reg net3 c_2_0 c_2_1 p_4 vdd1 vss1 full_adder
xi28 c_0_3_reg net22 c_1_2 c_1_3 s_1_3 vdd1 vss1 full_adder
xi22 s_0_3_reg net2 c_1_1 c_1_2 s_1_2 vdd1 vss1 full_adder
xi21 s_0_2_reg net4 c_1_0 c_1_1 s_1_1 vdd1 vss1 full_adder
xi14 net18 net35 c_0_1 c_0_2 s_0_2 vdd1 vss1 full_adder
xi13 net13 net45 c_0_0 c_0_1 s_0_1 vdd1 vss1 full_adder
xi125 p7_1_1 net59 vdd1 vss1 inverter_minsize
xi124 p3_1_1 net30 vdd1 vss1 inverter_minsize
xi123 p6_1_1 net53 vdd1 vss1 inverter_minsize
xi122 p2_1_1 net24 vdd1 vss1 inverter_minsize
xi121 p5_1_1 net47 vdd1 vss1 inverter_minsize
xi120 p1_1_1 net16 vdd1 vss1 inverter_minsize
xi119 p4_1_1 net38 vdd1 vss1 inverter_minsize
xi118 p0_1_1 net7 vdd1 vss1 inverter_minsize
xi90 clk_oc clk_bar vdd1 vss1 inverter_minsize
xi44 b_1_reg a_1_reg net45 vdd1 vss1 and_minsize
xi45 b_0_reg a_2_reg net13 vdd1 vss1 and_minsize
xi42 b_1_reg a_0_reg net8 vdd1 vss1 and_minsize
xi43 b_0_reg a_1_reg net10 vdd1 vss1 and_minsize
xi49 b_2_reg_reg a_0_reg_reg net5 vdd1 vss1 and_minsize
xi52 b_2_reg_reg a_3_reg_reg net22 vdd1 vss1 and_minsize
xi51 b_2_reg_reg a_2_reg_reg net2 vdd1 vss1 and_minsize
xi50 b_2_reg_reg a_1_reg_reg net4 vdd1 vss1 and_minsize
xi53 b_3_reg_reg_reg a_0_reg_reg_reg net6 vdd1 vss1 and_minsize
xi54 b_3_reg_reg_reg a_1_reg_reg_reg net3 vdd1 vss1 and_minsize
xi55 b_3_reg_reg_reg a_2_reg_reg_reg net1 vdd1 vss1 and_minsize
xi56 b_3_reg_reg_reg a_3_reg_reg_reg net11 vdd1 vss1 and_minsize
xi48 b_1_reg a_3_reg net41 vdd1 vss1 and_minsize
xi46 b_0_reg a_3_reg net18 vdd1 vss1 and_minsize
xi47 b_1_reg a_2_reg net35 vdd1 vss1 and_minsize
xi135 b_0_reg a_0_reg p_0 vdd1 vss1 and_minsize
xi75 rst_oc reset_bar rst rst_bar vdd1 vss1 level_shifter_1_8_to_1_1
xi74 b0_oc b0_bar b_0 b_0_bar vdd1 vss1 level_shifter_1_8_to_1_1
xi73 b1_oc b1_bar b_1 b_1_bar vdd1 vss1 level_shifter_1_8_to_1_1
xi72 b2_oc b2_bar b_2 b_2_bar vdd1 vss1 level_shifter_1_8_to_1_1
xi71 b3_oc b3_bar b_3 b_3_bar vdd1 vss1 level_shifter_1_8_to_1_1
xi70 a0_oc a0_bar a_0 a_0_bar vdd1 vss1 level_shifter_1_8_to_1_1
xi69 a1_oc a1_bar a_1 a_1_bar vdd1 vss1 level_shifter_1_8_to_1_1
xi68 a2_oc a2_bar a_2 a_2_bar vdd1 vss1 level_shifter_1_8_to_1_1
xi67 a3_oc a3_bar a_3 a_3_bar vdd1 vss1 level_shifter_1_8_to_1_1
xi84 rst_oc reset_bar vddio1 vss1 inverter_1_8_v
xi83 b0_oc b0_bar vddio1 vss1 inverter_1_8_v
xi82 b1_oc b1_bar vddio1 vss1 inverter_1_8_v
xi81 b2_oc b2_bar vddio1 vss1 inverter_1_8_v
xi80 b3_oc b3_bar vddio1 vss1 inverter_1_8_v
xi79 a0_oc a0_bar vddio1 vss1 inverter_1_8_v
xi78 a1_oc a1_bar vddio1 vss1 inverter_1_8_v
xi77 a2_oc a2_bar vddio1 vss1 inverter_1_8_v
xi76 a3_oc a3_bar vddio1 vss1 inverter_1_8_v
xi109 clk_oc clk_bar c_1_3 c_1_3_reg rst vdd1 vss1 C2MOS_register
xi108 clk_oc clk_bar s_1_3 s_1_3_reg rst vdd1 vss1 C2MOS_register
xi107 clk_oc clk_bar s_1_2 s_1_2_reg rst vdd1 vss1 C2MOS_register
xi106 clk_oc clk_bar s_1_1 s_1_1_reg rst vdd1 vss1 C2MOS_register
xi105 clk_oc clk_bar c_0_3 c_0_3_reg rst vdd1 vss1 C2MOS_register
xi104 clk_oc clk_bar s_0_3 s_0_3_reg rst vdd1 vss1 C2MOS_register
xi103 clk_oc clk_bar s_0_2 s_0_2_reg rst vdd1 vss1 C2MOS_register
xi102 clk_oc clk_bar s_0_1 s_0_1_reg rst vdd1 vss1 C2MOS_register
xi101 clk_oc clk_bar p_7 p7_1_1 rst vdd1 vss1 C2MOS_register
xi100 clk_oc clk_bar p_6 p6_1_1 rst vdd1 vss1 C2MOS_register
xi99 clk_oc clk_bar p_5 p5_1_1 rst vdd1 vss1 C2MOS_register
xi98 clk_oc clk_bar p_4 p4_1_1 rst vdd1 vss1 C2MOS_register
xi97 clk_oc clk_bar p_3 p3_1_1 rst vdd1 vss1 C2MOS_register
xi96 clk_oc clk_bar p_2 p_2_reg rst vdd1 vss1 C2MOS_register
xi95 clk_oc clk_bar p_2_reg p2_1_1 rst vdd1 vss1 C2MOS_register
xi94 clk_oc clk_bar p_1_reg p_1_reg_reg rst vdd1 vss1 C2MOS_register
xi93 clk_oc clk_bar p_0_reg p_0_reg_reg rst vdd1 vss1 C2MOS_register
xi92 clk_oc clk_bar p_1 p_1_reg rst vdd1 vss1 C2MOS_register
xi91 clk_oc clk_bar p_0 p_0_reg rst vdd1 vss1 C2MOS_register
xi89 clk_oc clk_bar a_3_reg_reg a_3_reg_reg_reg rst vdd1 vss1 C2MOS_register
xi88 clk_oc clk_bar a_2_reg_reg a_2_reg_reg_reg rst vdd1 vss1 C2MOS_register
xi87 clk_oc clk_bar a_1_reg_reg a_1_reg_reg_reg rst vdd1 vss1 C2MOS_register
xi86 clk_oc clk_bar a_0_reg_reg a_0_reg_reg_reg rst vdd1 vss1 C2MOS_register
xi85 clk_oc clk_bar b_3_reg_reg b_3_reg_reg_reg rst vdd1 vss1 C2MOS_register
xi66 clk_oc clk_bar b_3_reg b_3_reg_reg rst vdd1 vss1 C2MOS_register
xi65 clk_oc clk_bar b_2_reg b_2_reg_reg rst vdd1 vss1 C2MOS_register
xi64 clk_oc clk_bar a_3_reg a_3_reg_reg rst vdd1 vss1 C2MOS_register
xi63 clk_oc clk_bar a_2_reg a_2_reg_reg rst vdd1 vss1 C2MOS_register
xi60 clk_oc clk_bar p_1_reg_reg p1_1_1 rst vdd1 vss1 C2MOS_register
xi62 clk_oc clk_bar a_1_reg a_1_reg_reg rst vdd1 vss1 C2MOS_register
xi61 clk_oc clk_bar a_0_reg a_0_reg_reg rst vdd1 vss1 C2MOS_register
xi57 clk_oc clk_bar p_0_reg_reg p0_1_1 rst vdd1 vss1 C2MOS_register
xi7 clk_oc clk_bar b_3 b_3_reg rst vdd1 vss1 C2MOS_register
xi6 clk_oc clk_bar b_0 b_0_reg rst vdd1 vss1 C2MOS_register
xi5 clk_oc clk_bar b_1 b_1_reg rst vdd1 vss1 C2MOS_register
xi4 clk_oc clk_bar b_2 b_2_reg rst vdd1 vss1 C2MOS_register
xi3 clk_oc clk_bar a_0 a_0_reg rst vdd1 vss1 C2MOS_register
xi2 clk_oc clk_bar a_1 a_1_reg rst vdd1 vss1 C2MOS_register
xi1 clk_oc clk_bar a_2 a_2_reg rst vdd1 vss1 C2MOS_register
xi0 clk_oc clk_bar a_3 a_3_reg rst vdd1 vss1 C2MOS_register
xi160 vddio1 vss1 p7_f p7_oc superbuffer_4
xi158 vddio1 vss1 p2_f p2_oc superbuffer_4
xi155 vddio1 vss1 p4_f p4_oc superbuffer_4
xi154 vddio1 vss1 p0_f p0_oc superbuffer_4
xi159 vddio1 vss1 p6_f p6_oc superbuffer_4
xi156 vddio1 vss1 p5_f p5_oc superbuffer_4
xi157 vddio1 vss1 p1_f p1_oc superbuffer_4
xi161 vddio1 vss1 p3_f p3_oc superbuffer_4

*Put your extracted netlist above this comment













*Extracted PDN

** Library name: test2
** Cell name: pdn_rev3
** View name: av_extracted
xr41 rst_oc rst_oc1 resm11_pcell_0 segw=6e-6 segl=1e-6 dtemp=0
xr1 vdd2 vdd1 resm11_pcell_0 segw=6e-6 segl=1e-6 dtemp=0
xr0 vdd1 vdd2 resm11_pcell_0 segw=6e-6 segl=1e-6 dtemp=0
xr10 vddio1 vddio3 resm11_pcell_0 segw=6e-6 segl=1e-6 dtemp=0
xr11 vddio3 vddio1 resm11_pcell_0 segw=6e-6 segl=1e-6 dtemp=0
xr12 vss3 vss1 resm11_pcell_0 segw=6e-6 segl=1e-6 dtemp=0
xr13 vss1 vss3 resm11_pcell_0 segw=6e-6 segl=1e-6 dtemp=0
xr20 vss1 vssio3 resm11_pcell_0 segw=6e-6 segl=1e-6 dtemp=0
xr21 vssio3 vss1 resm11_pcell_0 segw=6e-6 segl=1e-6 dtemp=0
xr6 vdd1 vdd3 resm11_pcell_0 segw=6e-6 segl=1e-6 dtemp=0
xr7 vdd3 vdd1 resm11_pcell_0 segw=6e-6 segl=1e-6 dtemp=0
xr14 vss4 vss1 resm11_pcell_0 segw=6e-6 segl=1e-6 dtemp=0
xr15 vss1 vss4 resm11_pcell_0 segw=6e-6 segl=1e-6 dtemp=0
xr3 vddio2 vddio1 resm11_pcell_0 segw=6e-6 segl=1e-6 dtemp=0
xr2 vddio1 vddio2 resm11_pcell_0 segw=6e-6 segl=1e-6 dtemp=0
xr28 b0_oc b0_oc1 resm11_pcell_0 segw=6e-6 segl=1e-6 dtemp=0
xr29 b1_oc b1_oc1 resm11_pcell_0 segw=6e-6 segl=1e-6 dtemp=0
xr30 b2_oc b2_oc1 resm11_pcell_0 segw=6e-6 segl=1e-6 dtemp=0
xr31 b3_oc b3_oc1 resm11_pcell_0 segw=6e-6 segl=1e-6 dtemp=0
xr24 a0_oc a0_oc1 resm11_pcell_0 segw=6e-6 segl=1e-6 dtemp=0
xr25 a1_oc a1_oc1 resm11_pcell_0 segw=6e-6 segl=1e-6 dtemp=0
xr26 a2_oc a2_oc1 resm11_pcell_0 segw=6e-6 segl=1e-6 dtemp=0
xr27 a3_oc a3_oc1 resm11_pcell_0 segw=6e-6 segl=1e-6 dtemp=0
m80 _net0 _net1 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m81 _net0 _net1 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m82 _net2 _net3 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m83 _net2 _net3 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m84 _net8 _net9 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m85 _net8 _net9 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m86 _net10 _net11 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m87 _net10 _net11 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m88 _net10 _net11 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m89 _net8 _net9 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m90 _net10 _net11 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=450e-15 PD=6.4e-6 PS=6.3e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m91 _net8 _net9 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=450e-15 PD=6.4e-6 PS=6.3e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m92 _net2 _net3 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=450e-15 PD=6.4e-6 PS=6.3e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m93 _net0 _net1 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=450e-15 PD=6.4e-6 PS=6.3e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m94 _net2 _net3 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m95 _net0 _net1 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m96 _net4 _net5 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m97 _net4 _net5 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m98 _net6 _net7 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m99 _net6 _net7 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m100 _net12 _net13 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m101 _net12 _net13 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m102 _net14 _net15 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m103 _net14 _net15 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m104 _net14 _net15 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m105 _net12 _net13 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m106 _net14 _net15 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=450e-15 PD=6.4e-6 PS=6.3e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m107 _net12 _net13 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=450e-15 PD=6.4e-6 PS=6.3e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m108 _net6 _net7 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=450e-15 PD=6.4e-6 PS=6.3e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m109 _net4 _net5 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=450e-15 PD=6.4e-6 PS=6.3e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m110 _net6 _net7 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m111 _net4 _net5 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m112 _net16 _net17 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m113 _net16 _net17 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m114 _net18 _net19 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m115 _net18 _net19 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m116 _net24 _net25 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m117 _net24 _net25 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m118 _net26 _net27 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m119 _net26 _net27 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m120 _net26 _net27 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m121 _net24 _net25 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m122 _net26 _net27 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=450e-15 PD=6.4e-6 PS=6.3e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m123 _net24 _net25 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=450e-15 PD=6.4e-6 PS=6.3e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m124 _net18 _net19 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=450e-15 PD=6.4e-6 PS=6.3e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m125 _net16 _net17 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=450e-15 PD=6.4e-6 PS=6.3e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m126 _net18 _net19 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m127 _net16 _net17 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m128 _net20 _net21 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m129 _net20 _net21 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m130 _net22 _net23 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m131 _net22 _net23 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m132 _net28 _net29 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m133 _net28 _net29 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m134 _net30 _net31 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m135 _net30 _net31 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m136 _net30 _net31 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m137 _net28 _net29 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m138 _net30 _net31 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=450e-15 PD=6.4e-6 PS=6.3e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m139 _net28 _net29 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=450e-15 PD=6.4e-6 PS=6.3e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m140 _net22 _net23 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=450e-15 PD=6.4e-6 PS=6.3e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m141 _net20 _net21 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=450e-15 PD=6.4e-6 PS=6.3e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m142 _net22 _net23 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m143 _net20 _net21 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m144 _net32 _net33 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m145 _net32 _net33 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m146 _net34 _net35 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m147 _net34 _net35 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m148 _net40 _net41 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m149 _net40 _net41 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m150 _net42 _net43 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m151 _net42 _net43 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m152 _net42 _net43 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m153 _net40 _net41 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m154 _net42 _net43 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=450e-15 PD=6.4e-6 PS=6.3e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m155 _net40 _net41 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=450e-15 PD=6.4e-6 PS=6.3e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m156 _net34 _net35 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=450e-15 PD=6.4e-6 PS=6.3e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m157 _net32 _net33 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=450e-15 PD=6.4e-6 PS=6.3e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m158 _net34 _net35 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m159 _net32 _net33 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m160 _net36 _net37 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m161 _net36 _net37 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m162 _net38 _net39 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m163 _net38 _net39 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m164 _net44 _net45 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m165 _net44 _net45 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m166 _net46 _net47 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m167 _net46 _net47 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m168 _net46 _net47 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m169 _net44 _net45 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m170 _net46 _net47 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=450e-15 PD=6.4e-6 PS=6.3e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m171 _net44 _net45 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=450e-15 PD=6.4e-6 PS=6.3e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m172 _net38 _net39 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=450e-15 PD=6.4e-6 PS=6.3e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m173 _net36 _net37 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=450e-15 PD=6.4e-6 PS=6.3e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m174 _net38 _net39 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m175 _net36 _net37 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m176 _net48 _net49 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m177 _net48 _net49 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m178 _net50 _net51 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m179 _net50 _net51 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m180 _net56 _net57 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m181 _net56 _net57 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m182 _net58 _net59 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m183 _net58 _net59 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m184 _net58 _net59 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m185 _net56 _net57 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m186 _net58 _net59 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=450e-15 PD=6.4e-6 PS=6.3e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m187 _net56 _net57 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=450e-15 PD=6.4e-6 PS=6.3e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m188 _net50 _net51 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=450e-15 PD=6.4e-6 PS=6.3e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m189 _net48 _net49 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=450e-15 PD=6.4e-6 PS=6.3e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m190 _net50 _net51 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m191 _net48 _net49 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m192 _net52 _net53 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m193 _net52 _net53 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m194 _net54 _net55 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m195 _net54 _net55 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m196 _net60 _net61 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m197 _net60 _net61 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m198 _net62 _net63 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m199 _net62 _net63 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m200 _net62 _net63 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m201 _net60 _net61 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m202 _net62 _net63 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=450e-15 PD=6.4e-6 PS=6.3e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m203 _net60 _net61 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=450e-15 PD=6.4e-6 PS=6.3e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m204 _net54 _net55 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=450e-15 PD=6.4e-6 PS=6.3e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m205 _net52 _net53 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=450e-15 PD=6.4e-6 PS=6.3e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m206 _net54 _net55 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m207 _net52 _net53 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m208 _net64 _net65 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m209 _net64 _net65 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m210 _net66 _net67 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m211 _net66 _net67 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m212 _net72 _net73 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m213 _net72 _net73 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m214 _net74 _net75 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m215 _net74 _net75 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m216 _net74 _net75 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m217 _net72 _net73 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m218 _net74 _net75 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=450e-15 PD=6.4e-6 PS=6.3e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m219 _net72 _net73 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=450e-15 PD=6.4e-6 PS=6.3e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m220 _net66 _net67 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=450e-15 PD=6.4e-6 PS=6.3e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m221 _net64 _net65 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=450e-15 PD=6.4e-6 PS=6.3e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m222 _net66 _net67 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m223 _net64 _net65 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m224 _net68 _net69 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m225 _net68 _net69 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m226 _net70 _net71 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m227 _net70 _net71 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m228 _net76 _net77 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m229 _net76 _net77 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m230 _net78 _net79 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m231 _net78 _net79 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m232 _net78 _net79 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m233 _net76 _net77 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m234 _net78 _net79 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=450e-15 PD=6.4e-6 PS=6.3e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m235 _net76 _net77 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=450e-15 PD=6.4e-6 PS=6.3e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m236 _net70 _net71 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=450e-15 PD=6.4e-6 PS=6.3e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m237 _net68 _net69 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=450e-15 PD=6.4e-6 PS=6.3e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m238 _net70 _net71 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m239 _net68 _net69 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m240 _net78 _net79 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=450e-15 PD=6.4e-6 PS=6.3e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m241 _net76 _net77 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=450e-15 PD=6.4e-6 PS=6.3e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m242 _net74 _net75 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=450e-15 PD=6.4e-6 PS=6.3e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m243 _net72 _net73 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=450e-15 PD=6.4e-6 PS=6.3e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m244 _net78 _net79 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m245 _net76 _net77 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m246 _net74 _net75 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m247 _net72 _net73 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m248 _net70 _net71 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m249 _net68 _net69 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m250 _net66 _net67 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m251 _net64 _net65 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m252 _net70 _net71 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=450e-15 PD=6.4e-6 PS=6.3e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m253 _net68 _net69 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=450e-15 PD=6.4e-6 PS=6.3e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m254 _net66 _net67 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=450e-15 PD=6.4e-6 PS=6.3e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m255 _net64 _net65 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=450e-15 PD=6.4e-6 PS=6.3e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m256 _net62 _net63 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=450e-15 PD=6.4e-6 PS=6.3e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m257 _net60 _net61 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=450e-15 PD=6.4e-6 PS=6.3e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m258 _net58 _net59 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=450e-15 PD=6.4e-6 PS=6.3e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m259 _net56 _net57 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=450e-15 PD=6.4e-6 PS=6.3e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m260 _net62 _net63 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m261 _net60 _net61 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m262 _net58 _net59 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m263 _net56 _net57 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m264 _net54 _net55 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m265 _net52 _net53 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m266 _net50 _net51 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m267 _net48 _net49 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m268 _net54 _net55 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=450e-15 PD=6.4e-6 PS=6.3e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m269 _net52 _net53 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=450e-15 PD=6.4e-6 PS=6.3e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m270 _net50 _net51 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=450e-15 PD=6.4e-6 PS=6.3e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m271 _net48 _net49 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=450e-15 PD=6.4e-6 PS=6.3e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m272 _net46 _net47 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=450e-15 PD=6.4e-6 PS=6.3e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m273 _net44 _net45 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=450e-15 PD=6.4e-6 PS=6.3e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m274 _net42 _net43 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=450e-15 PD=6.4e-6 PS=6.3e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m275 _net40 _net41 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=450e-15 PD=6.4e-6 PS=6.3e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m276 _net46 _net47 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m277 _net44 _net45 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m278 _net42 _net43 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m279 _net40 _net41 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m280 _net38 _net39 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m281 _net36 _net37 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m282 _net34 _net35 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m283 _net32 _net33 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m284 _net38 _net39 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=450e-15 PD=6.4e-6 PS=6.3e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m285 _net36 _net37 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=450e-15 PD=6.4e-6 PS=6.3e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m286 _net34 _net35 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=450e-15 PD=6.4e-6 PS=6.3e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m287 _net32 _net33 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=450e-15 PD=6.4e-6 PS=6.3e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m288 _net30 _net31 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=450e-15 PD=6.4e-6 PS=6.3e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m289 _net28 _net29 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=450e-15 PD=6.4e-6 PS=6.3e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m290 _net26 _net27 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=450e-15 PD=6.4e-6 PS=6.3e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m291 _net24 _net25 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=450e-15 PD=6.4e-6 PS=6.3e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m292 _net30 _net31 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m293 _net28 _net29 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m294 _net26 _net27 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m295 _net24 _net25 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m296 _net22 _net23 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m297 _net20 _net21 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m298 _net18 _net19 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m299 _net16 _net17 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m300 _net22 _net23 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=450e-15 PD=6.4e-6 PS=6.3e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m301 _net20 _net21 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=450e-15 PD=6.4e-6 PS=6.3e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m302 _net18 _net19 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=450e-15 PD=6.4e-6 PS=6.3e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m303 _net16 _net17 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=450e-15 PD=6.4e-6 PS=6.3e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m304 _net14 _net15 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=450e-15 PD=6.4e-6 PS=6.3e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m305 _net12 _net13 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=450e-15 PD=6.4e-6 PS=6.3e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m306 _net10 _net11 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=450e-15 PD=6.4e-6 PS=6.3e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m307 _net8 _net9 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=450e-15 PD=6.4e-6 PS=6.3e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m308 _net14 _net15 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m309 _net12 _net13 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m310 _net10 _net11 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m311 _net8 _net9 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m312 _net6 _net7 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m313 _net4 _net5 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m314 _net2 _net3 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m315 _net0 _net1 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m316 _net6 _net7 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=450e-15 PD=6.4e-6 PS=6.3e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m317 _net4 _net5 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=450e-15 PD=6.4e-6 PS=6.3e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m318 _net2 _net3 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=450e-15 PD=6.4e-6 PS=6.3e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m319 _net0 _net1 vddio1 vddio1 g45p2svt L=150e-9 W=3e-6 AD=600e-15 AS=450e-15 PD=6.4e-6 PS=6.3e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
c1 a0_oc vss1 34.3825e-15
c2 a1_oc vss1 34.3825e-15
c3 a1_oc1 vss1 1.11514e-15
c4 a2_oc vss1 34.3825e-15
c5 a2_oc1 vss1 1.11514e-15
c6 a3_oc vss1 34.3825e-15
c7 a3_oc1 vss1 1.11514e-15
c8 a0_oc1 vss1 1.11514e-15
c9 b0_oc vss1 34.3825e-15
c10 b0_oc1 vss1 1.11514e-15
c11 b1_oc vss1 34.3825e-15
c12 b1_oc1 vss1 1.11514e-15
c13 b2_oc vss1 34.3825e-15
c14 b2_oc1 vss1 1.11514e-15
c15 b3_oc vss1 34.3825e-15
c16 b3_oc1 vss1 1.11514e-15
c17 clk_oc vss1 31.514e-15
c18 clk_oc1 vss1 1.43948e-15
c19 p0_oc vss1 33.9341e-15
c20 p0_oc1 vss1 1.3098e-15
c21 p1_oc vss1 33.9341e-15
c22 p1_oc1 vss1 1.3098e-15
c23 p2_oc vss1 33.9341e-15
c24 p2_oc1 vss1 1.3098e-15
c25 p3_oc vss1 33.9341e-15
c26 p3_oc1 vss1 1.3098e-15
c27 p4_oc vss1 33.9341e-15
c28 p4_oc1 vss1 1.3098e-15
c29 p5_oc vss1 33.9341e-15
c30 p5_oc1 vss1 1.3098e-15
c31 p6_oc vss1 33.9341e-15
c32 p6_oc1 vss1 1.3098e-15
c33 p7_oc vss1 33.9341e-15
c34 p7_oc1 vss1 1.3098e-15
c35 rst_oc vss1 34.3825e-15
c36 rst_oc1 vss1 1.11514e-15
c37 vdd1 vss1 70.8243e-12
c38 vdd2 vss1 835.125e-18
c39 vdd3 vss1 1.62092e-15
c40 vddio1 vss1 1.06771e-12
c41 vddio2 vss1 765.365e-18
c42 vddio3 vss1 1.15638e-15
c43 vss2 vss1 1.28488e-15
c44 vss3 vss1 907.659e-18
c45 vss4 vss1 1.03734e-15
c46 vssio1 vss1 1.15231e-15
c47 vssio2 vss1 1.36155e-15
c48 vssio3 vss1 1.16703e-15
c49 n16 vss1 32.6001e-15
c50 n18 vss1 32.6001e-15
c51 n20 vss1 32.6001e-15
c52 n22 vss1 32.6001e-15
c53 n24 vss1 32.6001e-15
c54 n26 vss1 32.6001e-15
c55 n28 vss1 29.4798e-15
c56 n29 vss1 29.4798e-15
c57 n30 vss1 29.4798e-15
c58 n31 vss1 29.4798e-15
c59 n32 vss1 29.4798e-15
c60 n33 vss1 29.4798e-15
c61 n34 vss1 29.4798e-15
c62 _net76 vss1 3.64447e-15
c63 _net78 vss1 3.59963e-15
c64 _net68 vss1 3.66559e-15
c65 _net70 vss1 3.61796e-15
c66 _net77 vss1 3.67553e-15
c67 _net79 vss1 3.7062e-15
c68 _net69 vss1 3.69324e-15
c69 _net71 vss1 3.72336e-15
c70 _net72 vss1 3.63875e-15
c71 _net74 vss1 3.59557e-15
c72 _net64 vss1 3.65668e-15
c73 _net66 vss1 3.61466e-15
c74 _net73 vss1 3.67559e-15
c75 _net75 vss1 3.70715e-15
c76 _net65 vss1 3.69247e-15
c77 _net67 vss1 3.72395e-15
c78 _net60 vss1 3.66253e-15
c79 _net62 vss1 3.61796e-15
c80 _net52 vss1 3.66253e-15
c81 _net54 vss1 3.61796e-15
c82 _net61 vss1 3.69269e-15
c83 _net63 vss1 3.72336e-15
c84 _net53 vss1 3.69269e-15
c85 _net55 vss1 3.72336e-15
c86 _net56 vss1 3.65667e-15
c87 _net58 vss1 3.61461e-15
c88 _net48 vss1 3.65673e-15
c89 _net50 vss1 3.61424e-15
c90 _net57 vss1 3.69213e-15
c91 _net59 vss1 3.72373e-15
c92 _net49 vss1 3.69226e-15
c93 _net51 vss1 3.72259e-15
c94 _net44 vss1 3.66688e-15
c95 _net46 vss1 3.61796e-15
c96 _net36 vss1 3.66272e-15
c97 _net38 vss1 3.61796e-15
c98 _net45 vss1 3.69398e-15
c99 _net47 vss1 3.72336e-15
c100 _net37 vss1 3.69269e-15
c101 _net39 vss1 3.72336e-15
c102 _net40 vss1 3.65693e-15
c103 _net42 vss1 3.61422e-15
c104 _net32 vss1 3.65667e-15
c105 _net34 vss1 3.61461e-15
c106 _net41 vss1 3.69223e-15
c107 _net43 vss1 3.7251e-15
c108 _net33 vss1 3.69213e-15
c109 _net35 vss1 3.72373e-15
c110 _net28 vss1 3.66253e-15
c111 _net30 vss1 3.61796e-15
c112 _net20 vss1 3.6648e-15
c113 _net22 vss1 3.61796e-15
c114 _net29 vss1 3.69269e-15
c115 _net31 vss1 3.72336e-15
c116 _net21 vss1 3.69401e-15
c117 _net23 vss1 3.72336e-15
c118 _net24 vss1 3.65667e-15
c119 _net26 vss1 3.61461e-15
c120 _net16 vss1 3.65698e-15
c121 _net18 vss1 3.61872e-15
c122 _net25 vss1 3.69215e-15
c123 _net27 vss1 3.72385e-15
c124 _net17 vss1 3.6923e-15
c125 _net19 vss1 3.72772e-15
c126 _net12 vss1 3.66226e-15
c127 _net14 vss1 3.61796e-15
c128 _net4 vss1 3.64421e-15
c129 _net6 vss1 3.59963e-15
c130 _net13 vss1 3.69269e-15
c131 _net15 vss1 3.72336e-15
c132 _net5 vss1 3.67765e-15
c133 _net7 vss1 3.70832e-15
c134 _net8 vss1 3.65667e-15
c135 _net10 vss1 3.61538e-15
c136 _net0 vss1 3.63834e-15
c137 _net2 vss1 3.59628e-15
c138 _net9 vss1 3.69213e-15
c139 _net11 vss1 3.72438e-15
c140 _net1 vss1 3.67709e-15
c141 _net3 vss1 3.7087e-15
m320 _net1 _net0 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=450e-15 PD=6.4e-6 PS=6.3e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m321 _net1 _net0 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m322 _net1 _net0 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m323 _net1 _net0 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m324 _net1 _net0 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m325 _net1 _net0 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=450e-15 PD=6.4e-6 PS=6.3e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m326 _net3 _net2 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=450e-15 PD=6.4e-6 PS=6.3e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m327 _net3 _net2 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m328 _net3 _net2 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m329 _net3 _net2 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m330 _net3 _net2 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m331 _net3 _net2 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=450e-15 PD=6.4e-6 PS=6.3e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m332 _net9 _net8 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=450e-15 PD=6.4e-6 PS=6.3e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m333 _net9 _net8 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m334 _net9 _net8 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m335 _net9 _net8 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m336 _net9 _net8 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m337 _net9 _net8 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=450e-15 PD=6.4e-6 PS=6.3e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m338 _net11 _net10 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=450e-15 PD=6.4e-6 PS=6.3e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m339 _net11 _net10 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m340 _net11 _net10 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m341 _net11 _net10 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m342 _net11 _net10 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m343 _net11 _net10 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=450e-15 PD=6.4e-6 PS=6.3e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m344 _net5 _net4 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=450e-15 PD=6.4e-6 PS=6.3e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m345 _net5 _net4 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m346 _net5 _net4 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m347 _net5 _net4 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m348 _net5 _net4 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m349 _net5 _net4 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=450e-15 PD=6.4e-6 PS=6.3e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m350 _net7 _net6 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=450e-15 PD=6.4e-6 PS=6.3e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m351 _net7 _net6 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m352 _net7 _net6 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m353 _net7 _net6 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m354 _net7 _net6 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m355 _net7 _net6 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=450e-15 PD=6.4e-6 PS=6.3e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m356 _net13 _net12 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=450e-15 PD=6.4e-6 PS=6.3e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m357 _net13 _net12 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m358 _net13 _net12 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m359 _net13 _net12 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m360 _net13 _net12 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m361 _net13 _net12 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=450e-15 PD=6.4e-6 PS=6.3e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m362 _net15 _net14 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=450e-15 PD=6.4e-6 PS=6.3e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m363 _net15 _net14 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m364 _net15 _net14 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m365 _net15 _net14 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m366 _net15 _net14 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m367 _net15 _net14 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=450e-15 PD=6.4e-6 PS=6.3e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m368 _net17 _net16 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=450e-15 PD=6.4e-6 PS=6.3e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m369 _net17 _net16 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m370 _net17 _net16 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m371 _net17 _net16 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m372 _net17 _net16 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m373 _net17 _net16 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=450e-15 PD=6.4e-6 PS=6.3e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m374 _net19 _net18 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=450e-15 PD=6.4e-6 PS=6.3e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m375 _net19 _net18 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m376 _net19 _net18 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m377 _net19 _net18 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m378 _net19 _net18 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m379 _net19 _net18 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=450e-15 PD=6.4e-6 PS=6.3e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m380 _net25 _net24 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=450e-15 PD=6.4e-6 PS=6.3e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m381 _net25 _net24 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m382 _net25 _net24 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m383 _net25 _net24 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m384 _net25 _net24 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m385 _net25 _net24 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=450e-15 PD=6.4e-6 PS=6.3e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m386 _net27 _net26 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=450e-15 PD=6.4e-6 PS=6.3e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m387 _net27 _net26 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m388 _net27 _net26 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m389 _net27 _net26 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m390 _net27 _net26 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m391 _net27 _net26 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=450e-15 PD=6.4e-6 PS=6.3e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m392 _net21 _net20 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=450e-15 PD=6.4e-6 PS=6.3e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m393 _net21 _net20 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m394 _net21 _net20 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m395 _net21 _net20 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m396 _net21 _net20 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m397 _net21 _net20 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=450e-15 PD=6.4e-6 PS=6.3e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m398 _net23 _net22 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=450e-15 PD=6.4e-6 PS=6.3e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m399 _net23 _net22 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m400 _net23 _net22 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m401 _net23 _net22 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m402 _net23 _net22 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m403 _net23 _net22 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=450e-15 PD=6.4e-6 PS=6.3e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m404 _net29 _net28 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=450e-15 PD=6.4e-6 PS=6.3e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m405 _net29 _net28 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m406 _net29 _net28 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m407 _net29 _net28 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m408 _net29 _net28 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m409 _net29 _net28 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=450e-15 PD=6.4e-6 PS=6.3e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m410 _net31 _net30 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=450e-15 PD=6.4e-6 PS=6.3e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m411 _net31 _net30 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m412 _net31 _net30 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m413 _net31 _net30 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m414 _net31 _net30 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m415 _net31 _net30 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=450e-15 PD=6.4e-6 PS=6.3e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m416 _net33 _net32 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=450e-15 PD=6.4e-6 PS=6.3e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m417 _net33 _net32 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m418 _net33 _net32 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m419 _net33 _net32 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m420 _net33 _net32 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m421 _net33 _net32 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=450e-15 PD=6.4e-6 PS=6.3e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m422 _net35 _net34 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=450e-15 PD=6.4e-6 PS=6.3e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m423 _net35 _net34 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m424 _net35 _net34 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m425 _net35 _net34 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m426 _net35 _net34 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m427 _net35 _net34 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=450e-15 PD=6.4e-6 PS=6.3e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m428 _net41 _net40 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=450e-15 PD=6.4e-6 PS=6.3e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m429 _net41 _net40 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m430 _net41 _net40 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m431 _net41 _net40 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m432 _net41 _net40 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m433 _net41 _net40 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=450e-15 PD=6.4e-6 PS=6.3e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m434 _net43 _net42 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=450e-15 PD=6.4e-6 PS=6.3e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m435 _net43 _net42 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m436 _net43 _net42 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m437 _net43 _net42 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m438 _net43 _net42 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m439 _net43 _net42 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=450e-15 PD=6.4e-6 PS=6.3e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m440 _net37 _net36 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=450e-15 PD=6.4e-6 PS=6.3e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m441 _net37 _net36 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m442 _net37 _net36 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m443 _net37 _net36 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m444 _net37 _net36 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m445 _net37 _net36 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=450e-15 PD=6.4e-6 PS=6.3e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m446 _net39 _net38 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=450e-15 PD=6.4e-6 PS=6.3e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m447 _net39 _net38 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m448 _net39 _net38 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m449 _net39 _net38 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m450 _net39 _net38 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m451 _net39 _net38 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=450e-15 PD=6.4e-6 PS=6.3e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m452 _net45 _net44 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=450e-15 PD=6.4e-6 PS=6.3e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m453 _net45 _net44 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m454 _net45 _net44 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m455 _net45 _net44 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m456 _net45 _net44 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m457 _net45 _net44 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=450e-15 PD=6.4e-6 PS=6.3e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m458 _net47 _net46 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=450e-15 PD=6.4e-6 PS=6.3e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m459 _net47 _net46 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m460 _net47 _net46 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m461 _net47 _net46 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m462 _net47 _net46 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m463 _net47 _net46 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=450e-15 PD=6.4e-6 PS=6.3e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m464 _net49 _net48 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=450e-15 PD=6.4e-6 PS=6.3e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m465 _net49 _net48 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m466 _net49 _net48 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m467 _net49 _net48 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m468 _net49 _net48 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m469 _net49 _net48 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=450e-15 PD=6.4e-6 PS=6.3e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m470 _net51 _net50 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=450e-15 PD=6.4e-6 PS=6.3e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m471 _net51 _net50 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m472 _net51 _net50 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m473 _net51 _net50 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m474 _net51 _net50 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m475 _net51 _net50 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=450e-15 PD=6.4e-6 PS=6.3e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m476 _net57 _net56 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=450e-15 PD=6.4e-6 PS=6.3e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m477 _net57 _net56 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m478 _net57 _net56 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m479 _net57 _net56 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m480 _net57 _net56 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m481 _net57 _net56 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=450e-15 PD=6.4e-6 PS=6.3e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m482 _net59 _net58 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=450e-15 PD=6.4e-6 PS=6.3e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m483 _net59 _net58 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m484 _net59 _net58 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m485 _net59 _net58 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m486 _net59 _net58 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m487 _net59 _net58 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=450e-15 PD=6.4e-6 PS=6.3e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m488 _net53 _net52 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=450e-15 PD=6.4e-6 PS=6.3e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m489 _net53 _net52 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m490 _net53 _net52 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m491 _net53 _net52 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m492 _net53 _net52 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m493 _net53 _net52 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=450e-15 PD=6.4e-6 PS=6.3e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m494 _net55 _net54 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=450e-15 PD=6.4e-6 PS=6.3e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m495 _net55 _net54 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m496 _net55 _net54 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m497 _net55 _net54 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m498 _net55 _net54 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m499 _net55 _net54 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=450e-15 PD=6.4e-6 PS=6.3e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m500 _net61 _net60 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=450e-15 PD=6.4e-6 PS=6.3e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m501 _net61 _net60 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m502 _net61 _net60 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m503 _net61 _net60 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m504 _net61 _net60 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m505 _net61 _net60 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=450e-15 PD=6.4e-6 PS=6.3e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m506 _net63 _net62 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=450e-15 PD=6.4e-6 PS=6.3e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m507 _net63 _net62 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m508 _net63 _net62 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m509 _net63 _net62 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m510 _net63 _net62 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m511 _net63 _net62 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=450e-15 PD=6.4e-6 PS=6.3e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m512 _net65 _net64 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=450e-15 PD=6.4e-6 PS=6.3e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m513 _net65 _net64 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m514 _net65 _net64 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m515 _net65 _net64 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m516 _net65 _net64 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m517 _net65 _net64 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=450e-15 PD=6.4e-6 PS=6.3e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m518 _net67 _net66 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=450e-15 PD=6.4e-6 PS=6.3e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m519 _net67 _net66 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m520 _net67 _net66 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m521 _net67 _net66 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m522 _net67 _net66 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m523 _net67 _net66 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=450e-15 PD=6.4e-6 PS=6.3e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m524 _net73 _net72 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=450e-15 PD=6.4e-6 PS=6.3e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m525 _net73 _net72 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m526 _net73 _net72 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m527 _net73 _net72 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m528 _net73 _net72 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m529 _net73 _net72 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=450e-15 PD=6.4e-6 PS=6.3e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m530 _net75 _net74 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=450e-15 PD=6.4e-6 PS=6.3e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m531 _net75 _net74 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m532 _net75 _net74 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m533 _net75 _net74 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m534 _net75 _net74 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m535 _net75 _net74 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=450e-15 PD=6.4e-6 PS=6.3e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m536 _net69 _net68 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=450e-15 PD=6.4e-6 PS=6.3e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m537 _net69 _net68 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m538 _net69 _net68 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m539 _net69 _net68 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m540 _net69 _net68 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m541 _net69 _net68 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=450e-15 PD=6.4e-6 PS=6.3e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m542 _net71 _net70 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=450e-15 PD=6.4e-6 PS=6.3e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m543 _net71 _net70 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m544 _net71 _net70 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m545 _net71 _net70 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m546 _net71 _net70 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m547 _net71 _net70 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=450e-15 PD=6.4e-6 PS=6.3e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m548 _net77 _net76 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=450e-15 PD=6.4e-6 PS=6.3e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m549 _net77 _net76 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m550 _net77 _net76 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m551 _net77 _net76 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m552 _net77 _net76 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m553 _net77 _net76 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=450e-15 PD=6.4e-6 PS=6.3e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m554 _net79 _net78 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=450e-15 PD=6.4e-6 PS=6.3e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m555 _net79 _net78 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m556 _net79 _net78 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m557 _net79 _net78 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m558 _net79 _net78 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=600e-15 PD=6.4e-6 PS=6.4e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
m559 _net79 _net78 vss1 vss1 g45n2svt L=150e-9 W=3e-6 AD=600e-15 AS=450e-15 PD=6.4e-6 PS=6.3e-6 NRD=468.75e-3 NRS=468.75e-3 M=1
xr5 vss1 vss2 resm11_pcell_0 segw=6e-6 segl=1e-6 dtemp=0
xr4 vss2 vss1 resm11_pcell_0 segw=6e-6 segl=1e-6 dtemp=0
xr39 p7_oc p7_oc1 resm11_pcell_0 segw=6e-6 segl=1e-6 dtemp=0
xr38 p6_oc p6_oc1 resm11_pcell_0 segw=6e-6 segl=1e-6 dtemp=0
xr37 p5_oc p5_oc1 resm11_pcell_0 segw=6e-6 segl=1e-6 dtemp=0
xr36 p4_oc p4_oc1 resm11_pcell_0 segw=6e-6 segl=1e-6 dtemp=0
xr35 p3_oc p3_oc1 resm11_pcell_0 segw=6e-6 segl=1e-6 dtemp=0
xr34 p2_oc p2_oc1 resm11_pcell_0 segw=6e-6 segl=1e-6 dtemp=0
xr33 p1_oc p1_oc1 resm11_pcell_0 segw=6e-6 segl=1e-6 dtemp=0
xr40 clk_oc clk_oc1 resm11_pcell_0 segw=6e-6 segl=1e-6 dtemp=0
xr32 p0_oc p0_oc1 resm11_pcell_0 segw=6e-6 segl=1e-6 dtemp=0
xr16 vss1 vssio1 resm11_pcell_0 segw=6e-6 segl=1e-6 dtemp=0
xr19 vss1 vssio2 resm11_pcell_0 segw=6e-6 segl=1e-6 dtemp=0
xr17 vssio1 vss1 resm11_pcell_0 segw=6e-6 segl=1e-6 dtemp=0
xr18 vssio2 vss1 resm11_pcell_0 segw=6e-6 segl=1e-6 dtemp=0





*End of Extracted PDN

* The load current required to be connected between the two terminals extracted from the netlist. You cannot modify it.
ILOAD vdd1 vss1 PWL(
+ 'tstart+0ns'      0mA    'tstart+0.25ns'   1.25mA   'tstart+0.5ns'    5mA     'tstart+0.75ns'   11.25mA
+ 'tstart+1ns'     20mA    'tstart+1.25ns'  28.75mA   'tstart+1.5ns'   35mA     'tstart+1.75ns'   38.75mA
+ 'tstart+2ns'     40mA    'tstart+2.25ns'  38.75mA   'tstart+2.5ns'   35mA     'tstart+2.75ns'   28.75mA
+ 'tstart+3ns'     20mA    'tstart+3.25ns'  11.25mA   'tstart+3.5ns'    5mA     'tstart+3.75ns'    1.25mA
+ 'tstart+4ns'      0mA    'tstart+4.25ns'   1.25mA   'tstart+4.5ns'    5mA     'tstart+4.75ns'   11.25mA
+ 'tstart+5ns'     20mA    'tstart+5.25ns'  28.75mA   'tstart+5.5ns'   35mA     'tstart+5.75ns'   38.75mA
+ 'tstart+6ns'     40mA    'tstart+6.25ns'  38.75mA   'tstart+6.5ns'   35mA     'tstart+6.75ns'   28.75mA
+ 'tstart+7ns'     20mA    'tstart+7.25ns'  11.25mA   'tstart+7.5ns'    5mA     'tstart+7.75ns'    1.25mA
+ 'tstart+8ns'      0mA    'tstart+8.25ns'   1.25mA   'tstart+8.5ns'    5mA     'tstart+8.75ns'   11.25mA
+ 'tstart+9ns'     20mA    'tstart+9.25ns'  28.75mA   'tstart+9.5ns'   35mA     'tstart+9.75ns'   38.75mA
+ 'tstart+10ns'    40mA    'tstart+10.25ns' 38.75mA   'tstart+10.5ns'  35mA     'tstart+10.75ns'  28.75mA
+ 'tstart+11ns'    20mA    'tstart+11.25ns' 11.25mA   'tstart+11.5ns'   5mA     'tstart+11.75ns'   1.25mA
+ 'tstart+12ns'     0mA    'tstart+12.25ns'  1.25mA   'tstart+12.5ns'   5mA     'tstart+12.75ns'  11.25mA
+ 'tstart+13ns'    20mA    'tstart+13.25ns' 28.75mA   'tstart+13.5ns'  35mA     'tstart+13.75ns'  38.75mA
+ 'tstart+14ns'    40mA    'tstart+14.25ns' 38.75mA   'tstart+14.5ns'  35mA     'tstart+14.75ns'  28.75mA
+ 'tstart+15ns'    20mA    'tstart+15.25ns' 11.25mA   'tstart+15.5ns'   5mA     'tstart+15.75ns'   1.25mA
+ 'tstart+16ns'     0mA    'tstart+16.25ns'  1.25mA   'tstart+16.5ns'   5mA     'tstart+16.75ns'  11.25mA
+ 'tstart+17ns'    20mA    'tstart+17.25ns' 28.75mA   'tstart+17.5ns'  35mA     'tstart+17.75ns'  38.75mA
+ 'tstart+18ns'    40mA    'tstart+18.25ns' 38.75mA   'tstart+18.5ns'  35mA     'tstart+18.75ns'  28.75mA
+ 'tstart+19ns'    20mA    'tstart+19.25ns' 11.25mA   'tstart+19.5ns'   5mA     'tstart+19.75ns'   1.25mA
+ 'tstart+20ns'     0mA    'tstart+20.25ns'  1.25mA   'tstart+20.5ns'   5mA     'tstart+20.75ns'  11.25mA
+ 'tstart+21ns'    20mA    'tstart+21.25ns' 28.75mA   'tstart+21.5ns'  35mA     'tstart+21.75ns'  38.75mA
+ 'tstart+22ns'    40mA    'tstart+22.25ns' 38.75mA   'tstart+22.5ns'  35mA     'tstart+22.75ns'  28.75mA
+ 'tstart+23ns'    20mA    'tstart+23.25ns' 11.25mA   'tstart+23.5ns'   5mA     'tstart+23.75ns'   1.25mA
+ 'tstart+24ns'     0mA    'tstart+24.25ns'  1.25mA   'tstart+24.5ns'   5mA     'tstart+24.75ns'  11.25mA
+ 'tstart+25ns'    20mA    'tstart+25.25ns' 28.75mA   'tstart+25.5ns'  35mA     'tstart+25.75ns'  38.75mA
+ 'tstart+26ns'    40mA    'tstart+26.25ns' 38.75mA   'tstart+26.5ns'  35mA     'tstart+26.75ns'  28.75mA
+ 'tstart+27ns'    20mA    'tstart+27.25ns' 11.25mA   'tstart+27.5ns'   5mA     'tstart+27.75ns'   1.25mA
+ 'tstart+28ns'     0mA    'tstart+28.25ns'  1.25mA   'tstart+28.5ns'   5mA     'tstart+28.75ns'  11.25mA
+ 'tstart+29ns'    20mA    'tstart+29.25ns' 28.75mA   'tstart+29.5ns'  35mA     'tstart+29.75ns'  38.75mA
+ 'tstart+30ns'    40mA    'tstart+30.25ns' 38.75mA   'tstart+30.5ns'  35mA     'tstart+30.75ns'  28.75mA
+ 'tstart+31ns'    20mA    'tstart+31.25ns' 11.25mA   'tstart+31.5ns'   5mA     'tstart+31.75ns'   1.25mA
+ 'tstart+32ns'     0mA    'tstart+32.25ns'  1.25mA   'tstart+32.5ns'   5mA     'tstart+32.75ns'  11.25mA
+ 'tstart+33ns'    20mA    'tstart+33.25ns' 28.75mA   'tstart+33.5ns'  35mA     'tstart+33.75ns'  38.75mA
+ 'tstart+34ns'    40mA    'tstart+34.25ns' 38.75mA   'tstart+34.5ns'  35mA     'tstart+34.75ns'  28.75mA
+ 'tstart+35ns'    20mA    'tstart+35.25ns' 11.25mA   'tstart+35.5ns'   5mA     'tstart+35.75ns'   1.25mA
+ 'tstart+36ns'     0mA    'tstart+36.25ns'  1.25mA   'tstart+36.5ns'   5mA     'tstart+36.75ns'  11.25mA
+ 'tstart+37ns'    20mA    'tstart+37.25ns' 28.75mA   'tstart+37.5ns'  35mA     'tstart+37.75ns'  38.75mA
+ 'tstart+38ns'    40mA    'tstart+38.25ns' 38.75mA   'tstart+38.5ns'  35mA     'tstart+38.75ns'  28.75mA
+ 'tstart+39ns'    20mA    'tstart+39.25ns' 11.25mA   'tstart+39.5ns'   5mA     'tstart+39.75ns'   1.25mA
+ 'tstart+40ns'     0mA
)



*Clock and reset signal
vCK clk_in 0 pulse(0 1.1 trf_ck trf_ck trf_ck CK_pw TCK)
vReset reset 0 PWL(0 1.8 reset_delay 1.8 'reset_delay+trf_ip_reset' 1.8 'reset_delay+reset_pw+trf_ip_reset' 1.8 'reset_delay+reset_pw+2*trf_ip_reset' 0 'reset_delay+reset_pw+2*trf_ip_reset+reset_delay2' 0 'reset_delay+reset_pw+3*trf_ip_reset+reset_delay2' 1.8 'reset_delay+2*reset_pw+3*trf_ip_reset+reset_delay2' 1.8 'reset_delay+2*reset_pw+4*trf_ip_reset+reset_delay2' 0 sim_end 0)

*Clock buffer
mnm1 clk net31782 vss vss g45n1svt L=45e-9 W=9.6e-6 AD=768e-15 AS=825.6e-15 PD=12.8e-6 PS=14e-6 NRD=8.33333e-3 NRS=8.95833e-3 M=1
mnm0 net31782 clk_in vss vss g45n1svt L=45e-9 W=2.4e-6 AD=192e-15 AS=206.4e-15 PD=5.6e-6 PS=6.08e-6 NRD=33.3333e-3 NRS=35.8333e-3 M=1
mpm1 clk net31782 vdd vdd g45p1svt L=45e-9 W=19.2e-6 AD=1.536e-12 AS=1.6512e-12 PD=22.4e-6 PS=24.56e-6 NRD=4.16667e-3 NRS=4.47917e-3 M=1
mpm0 net31782 clk_in vdd vdd g45p1svt L=45e-9 W=4.8e-6 AD=384e-15 AS=412.8e-15 PD=8e-6 PS=8.72e-6 NRD=16.6667e-3 NRS=17.9167e-3 M=1

*Input signals
vA2 a2 0 PWL(0 0 'input_delay+0*trf_ip_reset+0*input_pw' 0 'input_delay+1*trf_ip_reset+0*input_pw' 1.8 'input_delay+1*trf_ip_reset+1*input_pw' 1.8 'input_delay+2*trf_ip_reset+1*input_pw' 0 'input_delay+2*trf_ip_reset+2*input_pw' 0 'input_delay+3*trf_ip_reset+2*input_pw' 1.8 'input_delay+3*trf_ip_reset+3*input_pw' 1.8  'input_delay+4*trf_ip_reset+3*input_pw' 1.8 'input_delay+4*trf_ip_reset+4*input_pw' 1.8 'input_delay+5*trf_ip_reset+4*input_pw' 0 sim_end 0)
vA0 a0 0 PWL(0 0 'input_delay2+0*trf_ip_reset+0*input_pw' 0 'input_delay2+1*trf_ip_reset+0*input_pw' 1.8 'input_delay2+1*trf_ip_reset+1*input_pw' 1.8 'input_delay2+2*trf_ip_reset+1*input_pw' 1.8 'input_delay2+2*trf_ip_reset+2*input_pw' 1.8 'input_delay2+3*trf_ip_reset+2*input_pw' 1.8 'input_delay2+3*trf_ip_reset+3*input_pw' 1.8  'input_delay2+4*trf_ip_reset+3*input_pw' 0 'input_delay2+4*trf_ip_reset+4*input_pw' 0 'input_delay2+5*trf_ip_reset+4*input_pw' 1.8 sim_end 1.8)
vA3 a3 0 PWL(0 0 'input_delay3+0*trf_ip_reset+0*input_pw' 0 'input_delay3+1*trf_ip_reset+0*input_pw' 0 'input_delay3+1*trf_ip_reset+1*input_pw' 0 'input_delay3+2*trf_ip_reset+1*input_pw' 0 'input_delay3+2*trf_ip_reset+2*input_pw' 0 'input_delay3+3*trf_ip_reset+2*input_pw' 1.8 'input_delay3+3*trf_ip_reset+3*input_pw' 1.8  'input_delay3+4*trf_ip_reset+3*input_pw' 0 'input_delay3+4*trf_ip_reset+4*input_pw' 0 'input_delay3+5*trf_ip_reset+4*input_pw' 1.8 sim_end 1.8)
vA1 a1 0 PWL(0 0 'input_delay4+0*trf_ip_reset+0*input_pw' 0 'input_delay4+1*trf_ip_reset+0*input_pw' 1.8 'input_delay4+1*trf_ip_reset+1*input_pw' 1.8 'input_delay4+2*trf_ip_reset+1*input_pw' 1.8 'input_delay4+2*trf_ip_reset+2*input_pw' 1.8 'input_delay4+3*trf_ip_reset+2*input_pw' 1.8 'input_delay4+3*trf_ip_reset+3*input_pw' 1.8  'input_delay4+4*trf_ip_reset+3*input_pw' 1.8 'input_delay4+4*trf_ip_reset+4*input_pw' 1.8 'input_delay4+5*trf_ip_reset+4*input_pw' 0 sim_end 0)
vB3 b3 0 PWL(0 0 'input_delay2+0*trf_ip_reset+0*input_pw' 0 'input_delay2+1*trf_ip_reset+0*input_pw' 1.8 'input_delay2+1*trf_ip_reset+1*input_pw' 1.8 'input_delay2+2*trf_ip_reset+1*input_pw' 1.8 'input_delay2+2*trf_ip_reset+2*input_pw' 1.8 'input_delay2+3*trf_ip_reset+2*input_pw' 1.8 'input_delay2+3*trf_ip_reset+3*input_pw' 1.8  'input_delay2+4*trf_ip_reset+3*input_pw' 0 'input_delay2+4*trf_ip_reset+4*input_pw' 0 'input_delay2+5*trf_ip_reset+4*input_pw' 1.8 sim_end 1.8)
vB1 b1 0 PWL(0 0 'input_delay+0*trf_ip_reset+0*input_pw' 0 'input_delay+1*trf_ip_reset+0*input_pw' 0 'input_delay+1*trf_ip_reset+1*input_pw' 0 'input_delay+2*trf_ip_reset+1*input_pw' 0 'input_delay+2*trf_ip_reset+2*input_pw' 0 'input_delay+2*trf_ip_reset+2*input_pw+offset_ip' 0 'input_delay+3*trf_ip_reset+2*input_pw+offset_ip' 1.8 'input_delay+3*trf_ip_reset+3*input_pw+offset_ip' 1.8  'input_delay+4*trf_ip_reset+3*input_pw+offset_ip' 1.8 'input_delay+4*trf_ip_reset+4*input_pw+offset_ip' 1.8 'input_delay+5*trf_ip_reset+4*input_pw+offset_ip' 1.8 sim_end 1.8)
vB0 b0 0 PWL(0 0 'input_delay2+0*trf_ip_reset+0*input_pw' 0 'input_delay2+1*trf_ip_reset+0*input_pw' 0 'input_delay2+1*trf_ip_reset+1*input_pw' 0 'input_delay2+2*trf_ip_reset+1*input_pw' 1.8 'input_delay2+2*trf_ip_reset+2*input_pw' 1.8 'input_delay2+3*trf_ip_reset+2*input_pw' 1.8 'input_delay2+3*trf_ip_reset+3*input_pw' 1.8  'input_delay2+4*trf_ip_reset+3*input_pw' 0 'input_delay2+4*trf_ip_reset+4*input_pw' 0 'input_delay2+5*trf_ip_reset+4*input_pw' 1.8 sim_end 1.8)
vB2 b2 0 PWL(0 0 'input_delay4+0*trf_ip_reset+0*input_pw' 0 'input_delay4+1*trf_ip_reset+0*input_pw' 0 'input_delay4+1*trf_ip_reset+1*input_pw' 0 'input_delay4+2*trf_ip_reset+1*input_pw' 0 'input_delay4+2*trf_ip_reset+2*input_pw' 0 'input_delay4+3*trf_ip_reset+2*input_pw' 1.8 'input_delay4+3*trf_ip_reset+3*input_pw' 1.8  'input_delay4+4*trf_ip_reset+3*input_pw' 1.8 'input_delay4+4*trf_ip_reset+4*input_pw' 1.8 'input_delay4+5*trf_ip_reset+4*input_pw' 1.8 sim_end 1.8)

*Sources on board - ONly nom_vdd value can be modified for power reduction using the parameters above.
vVDDIO VDDIO 0 1.8
vVDD VDD 0 nom_vdd
vVSS VSS 0 0

*Bondwire inductance - Not to be modified.
LVSS1 vss1 VSS 2.5n
LVSS2 vss2 VSS 2.5n
LVSS3 vss3 VSS 2.5n
LVSS4 vss4 VSS 2.5n
LVSSIO1 vssio1 VSS 2.5n
LVSSIO2 vssio2 VSS 2.5n
LVSSIO3 vssio3 VSS 2.5n
LVDDIO1 vddio1 VDDIO 5n
LVDDIO2 vddio2 VDDIO 5n
LVDDIO3 vddio3 VDDIO 5n
LVDD1 vdd1 VDD 5n
LVDD2 vdd2 VDD 5n
LVDD3 vdd3 VDD 5n

LA0 a0 a0_oc 4n
LA1 a1 a1_oc 4n
LA2 a2 a2_oc 4n
LA3 a3 a3_oc 4n
LB0 b0 b0_oc 4n
LB1 b1 b1_oc 4n
LB2 b2 b2_oc 4n
LB3 b3 b3_oc 4n

LP0 p0 p0_oc 4n
LP1 p1 p1_oc 4n
LP2 p2 p2_oc 4n
LP3 p3 p3_oc 4n
LP4 p4 p4_oc 4n
LP5 p5 p5_oc 4n
LP6 p6 p6_oc 4n
LP7 p7 p7_oc 4n

LRST reset rst_oc 4n
LCLK clk clk_oc 2n

*ESD capacitance - Not to be modified.
CVDD1 vdd1 vss1 0.3p
CVDD2 vdd2 vss2 0.3p
CVDD3 vdd3 vss3 0.3p
CVDDIO1 vdd1 vss1 0.4p
CVDDIO2 vdd2 vss2 0.4p
CVDDIO3 vdd3 vss3 0.4p

CA0_OC a0_oc1 vss4 0.25p
CA1_OC a1_oc1 vssio1 0.25p
CA2_OC a2_oc1 vssio2 0.25p
CA3_OC a3_oc1 vssio3 0.25p
CB0_OC b0_oc1 vss1 0.25p
CB1_OC b1_oc1 vss2 0.25p
CB2_OC b2_oc1 vss3 0.25p
CB3_OC b3_oc1 vss4 0.25p

CP0_OC p0_oc1 vss4 0.25p
CP1_OC p1_oc1 vssio1 0.25p
CP2_OC p2_oc1 vssio2 0.25p
CP3_OC p3_oc1 vssio3 0.25p
CP4_OC p4_oc1 vss1 0.25p
CP5_OC p5_oc1 vss2 0.25p
CP6_OC p6_oc1 vss3 0.25p
CP7_OC p7_oc1 vss4 0.25p


CCLK_OC clk_oc1 vss1 0.3p
CRST_OC rst_oc1 vss1 0.25p

*Load Capacitance - Not to be modified.
CA0 a0 VSS 20p
CA1 a1 VSS 20p
CA2 a2 VSS 20p
CA3 a3 VSS 20p
CB0 b0 VSS 20p
CB1 b1 VSS 20p
CB2 b2 VSS 20p
CB3 b3 VSS 20p

CP0 p0 VSS 20p
CP1 p1 VSS 20p
CP2 p2 VSS 20p
CP3 p3 VSS 20p
CP4 p4 VSS 20p
CP5 p5 VSS 20p
CP6 p6 VSS 20p
CP7 p7 VSS 20p


CCLK clk VSS 2p
CRST reset VSS 20p

.tran 0 sim_end

*Power measurement functions - NOt to be modified.
.meas tran avg_pwr_vdd avg p(vVDD) from=reset_delay+reset_pw+2*trf_ip_reset to=sim_end-2n
.meas tran avg_pwr_vddio avg p(vVDDIO) from=reset_delay+reset_pw+2*trf_ip_reset to=sim_end-2n
* Corrected power after subtracting noisy current source power
.meas tran corrected_pwr_vdd  param='avg_pwr_vdd + 0.0217681251338'

.probe tran i(ILOAD)
.print tran vdd_net='v(vdd1) - v(vss1)'
.print tran vddio_net='v(vddio1) - v(vssio1)'
.option post
.end
