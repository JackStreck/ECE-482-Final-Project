ECE 482 PROJECT TESTBENCH
.lib '/class/ece482/gpdk045_mos' TT
.include "resm11_pcell_1.sp"

*The following parameter can be modified.
.param nom_vdd = 1.1

*The following parameters cannot be modified.
.param tstart = 1n
.param TCK = 4n
.param trf_ck = 200p
.param trf_ip_reset = 200p
.param reset_pw = 6n
.param CK_pw = 0.5*TCK
.param reset_delay = 1n
.param reset_delay2 = 10n
.param sim_end = 11*TCK
.param input_delay = 9.5n
.param input_delay2 = 9.7n
.param input_delay3 = 9.2n
.param input_delay4 = 9.8n
.param input_pw = 1*TCK
.param offset_ip = 1n

*Put your extracted netlist below this comment

*Put your extracted netlist above this comment

* The load current required to be connected between the two terminals extracted from the netlist. You cannot modify it.
ILOAD vdd1 vss1 PWL(
+ 'tstart+0ns'      0mA    'tstart+0.25ns'   1.25mA   'tstart+0.5ns'    5mA     'tstart+0.75ns'   11.25mA
+ 'tstart+1ns'     20mA    'tstart+1.25ns'  28.75mA   'tstart+1.5ns'   35mA     'tstart+1.75ns'   38.75mA
+ 'tstart+2ns'     40mA    'tstart+2.25ns'  38.75mA   'tstart+2.5ns'   35mA     'tstart+2.75ns'   28.75mA
+ 'tstart+3ns'     20mA    'tstart+3.25ns'  11.25mA   'tstart+3.5ns'    5mA     'tstart+3.75ns'    1.25mA
+ 'tstart+4ns'      0mA    'tstart+4.25ns'   1.25mA   'tstart+4.5ns'    5mA     'tstart+4.75ns'   11.25mA
+ 'tstart+5ns'     20mA    'tstart+5.25ns'  28.75mA   'tstart+5.5ns'   35mA     'tstart+5.75ns'   38.75mA
+ 'tstart+6ns'     40mA    'tstart+6.25ns'  38.75mA   'tstart+6.5ns'   35mA     'tstart+6.75ns'   28.75mA
+ 'tstart+7ns'     20mA    'tstart+7.25ns'  11.25mA   'tstart+7.5ns'    5mA     'tstart+7.75ns'    1.25mA
+ 'tstart+8ns'      0mA    'tstart+8.25ns'   1.25mA   'tstart+8.5ns'    5mA     'tstart+8.75ns'   11.25mA
+ 'tstart+9ns'     20mA    'tstart+9.25ns'  28.75mA   'tstart+9.5ns'   35mA     'tstart+9.75ns'   38.75mA
+ 'tstart+10ns'    40mA    'tstart+10.25ns' 38.75mA   'tstart+10.5ns'  35mA     'tstart+10.75ns'  28.75mA
+ 'tstart+11ns'    20mA    'tstart+11.25ns' 11.25mA   'tstart+11.5ns'   5mA     'tstart+11.75ns'   1.25mA
+ 'tstart+12ns'     0mA    'tstart+12.25ns'  1.25mA   'tstart+12.5ns'   5mA     'tstart+12.75ns'  11.25mA
+ 'tstart+13ns'    20mA    'tstart+13.25ns' 28.75mA   'tstart+13.5ns'  35mA     'tstart+13.75ns'  38.75mA
+ 'tstart+14ns'    40mA    'tstart+14.25ns' 38.75mA   'tstart+14.5ns'  35mA     'tstart+14.75ns'  28.75mA
+ 'tstart+15ns'    20mA    'tstart+15.25ns' 11.25mA   'tstart+15.5ns'   5mA     'tstart+15.75ns'   1.25mA
+ 'tstart+16ns'     0mA    'tstart+16.25ns'  1.25mA   'tstart+16.5ns'   5mA     'tstart+16.75ns'  11.25mA
+ 'tstart+17ns'    20mA    'tstart+17.25ns' 28.75mA   'tstart+17.5ns'  35mA     'tstart+17.75ns'  38.75mA
+ 'tstart+18ns'    40mA    'tstart+18.25ns' 38.75mA   'tstart+18.5ns'  35mA     'tstart+18.75ns'  28.75mA
+ 'tstart+19ns'    20mA    'tstart+19.25ns' 11.25mA   'tstart+19.5ns'   5mA     'tstart+19.75ns'   1.25mA
+ 'tstart+20ns'     0mA    'tstart+20.25ns'  1.25mA   'tstart+20.5ns'   5mA     'tstart+20.75ns'  11.25mA
+ 'tstart+21ns'    20mA    'tstart+21.25ns' 28.75mA   'tstart+21.5ns'  35mA     'tstart+21.75ns'  38.75mA
+ 'tstart+22ns'    40mA    'tstart+22.25ns' 38.75mA   'tstart+22.5ns'  35mA     'tstart+22.75ns'  28.75mA
+ 'tstart+23ns'    20mA    'tstart+23.25ns' 11.25mA   'tstart+23.5ns'   5mA     'tstart+23.75ns'   1.25mA
+ 'tstart+24ns'     0mA    'tstart+24.25ns'  1.25mA   'tstart+24.5ns'   5mA     'tstart+24.75ns'  11.25mA
+ 'tstart+25ns'    20mA    'tstart+25.25ns' 28.75mA   'tstart+25.5ns'  35mA     'tstart+25.75ns'  38.75mA
+ 'tstart+26ns'    40mA    'tstart+26.25ns' 38.75mA   'tstart+26.5ns'  35mA     'tstart+26.75ns'  28.75mA
+ 'tstart+27ns'    20mA    'tstart+27.25ns' 11.25mA   'tstart+27.5ns'   5mA     'tstart+27.75ns'   1.25mA
+ 'tstart+28ns'     0mA    'tstart+28.25ns'  1.25mA   'tstart+28.5ns'   5mA     'tstart+28.75ns'  11.25mA
+ 'tstart+29ns'    20mA    'tstart+29.25ns' 28.75mA   'tstart+29.5ns'  35mA     'tstart+29.75ns'  38.75mA
+ 'tstart+30ns'    40mA    'tstart+30.25ns' 38.75mA   'tstart+30.5ns'  35mA     'tstart+30.75ns'  28.75mA
+ 'tstart+31ns'    20mA    'tstart+31.25ns' 11.25mA   'tstart+31.5ns'   5mA     'tstart+31.75ns'   1.25mA
+ 'tstart+32ns'     0mA    'tstart+32.25ns'  1.25mA   'tstart+32.5ns'   5mA     'tstart+32.75ns'  11.25mA
+ 'tstart+33ns'    20mA    'tstart+33.25ns' 28.75mA   'tstart+33.5ns'  35mA     'tstart+33.75ns'  38.75mA
+ 'tstart+34ns'    40mA    'tstart+34.25ns' 38.75mA   'tstart+34.5ns'  35mA     'tstart+34.75ns'  28.75mA
+ 'tstart+35ns'    20mA    'tstart+35.25ns' 11.25mA   'tstart+35.5ns'   5mA     'tstart+35.75ns'   1.25mA
+ 'tstart+36ns'     0mA    'tstart+36.25ns'  1.25mA   'tstart+36.5ns'   5mA     'tstart+36.75ns'  11.25mA
+ 'tstart+37ns'    20mA    'tstart+37.25ns' 28.75mA   'tstart+37.5ns'  35mA     'tstart+37.75ns'  38.75mA
+ 'tstart+38ns'    40mA    'tstart+38.25ns' 38.75mA   'tstart+38.5ns'  35mA     'tstart+38.75ns'  28.75mA
+ 'tstart+39ns'    20mA    'tstart+39.25ns' 11.25mA   'tstart+39.5ns'   5mA     'tstart+39.75ns'   1.25mA
+ 'tstart+40ns'     0mA
)



*Clock and reset signal
vCK clk_in 0 pulse(0 1.1 trf_ck trf_ck trf_ck CK_pw TCK)
vReset reset 0 PWL(0 1.8 reset_delay 1.8 'reset_delay+trf_ip_reset' 1.8 'reset_delay+reset_pw+trf_ip_reset' 1.8 'reset_delay+reset_pw+2*trf_ip_reset' 0 'reset_delay+reset_pw+2*trf_ip_reset+reset_delay2' 0 'reset_delay+reset_pw+3*trf_ip_reset+reset_delay2' 1.8 'reset_delay+2*reset_pw+3*trf_ip_reset+reset_delay2' 1.8 'reset_delay+2*reset_pw+4*trf_ip_reset+reset_delay2' 0 sim_end 0)

*Clock buffer
mnm1 clk net31782 vss vss g45n1svt L=45e-9 W=9.6e-6 AD=768e-15 AS=825.6e-15 PD=12.8e-6 PS=14e-6 NRD=8.33333e-3 NRS=8.95833e-3 M=1
mnm0 net31782 clk_in vss vss g45n1svt L=45e-9 W=2.4e-6 AD=192e-15 AS=206.4e-15 PD=5.6e-6 PS=6.08e-6 NRD=33.3333e-3 NRS=35.8333e-3 M=1
mpm1 clk net31782 vdd vdd g45p1svt L=45e-9 W=19.2e-6 AD=1.536e-12 AS=1.6512e-12 PD=22.4e-6 PS=24.56e-6 NRD=4.16667e-3 NRS=4.47917e-3 M=1
mpm0 net31782 clk_in vdd vdd g45p1svt L=45e-9 W=4.8e-6 AD=384e-15 AS=412.8e-15 PD=8e-6 PS=8.72e-6 NRD=16.6667e-3 NRS=17.9167e-3 M=1

*Input signals
vA2 a2 0 PWL(0 0 'input_delay+0*trf_ip_reset+0*input_pw' 0 'input_delay+1*trf_ip_reset+0*input_pw' 1.8 'input_delay+1*trf_ip_reset+1*input_pw' 1.8 'input_delay+2*trf_ip_reset+1*input_pw' 0 'input_delay+2*trf_ip_reset+2*input_pw' 0 'input_delay+3*trf_ip_reset+2*input_pw' 1.8 'input_delay+3*trf_ip_reset+3*input_pw' 1.8  'input_delay+4*trf_ip_reset+3*input_pw' 1.8 'input_delay+4*trf_ip_reset+4*input_pw' 1.8 'input_delay+5*trf_ip_reset+4*input_pw' 0 sim_end 0)
vA0 a0 0 PWL(0 0 'input_delay2+0*trf_ip_reset+0*input_pw' 0 'input_delay2+1*trf_ip_reset+0*input_pw' 1.8 'input_delay2+1*trf_ip_reset+1*input_pw' 1.8 'input_delay2+2*trf_ip_reset+1*input_pw' 1.8 'input_delay2+2*trf_ip_reset+2*input_pw' 1.8 'input_delay2+3*trf_ip_reset+2*input_pw' 1.8 'input_delay2+3*trf_ip_reset+3*input_pw' 1.8  'input_delay2+4*trf_ip_reset+3*input_pw' 0 'input_delay2+4*trf_ip_reset+4*input_pw' 0 'input_delay2+5*trf_ip_reset+4*input_pw' 1.8 sim_end 1.8)
vA3 a3 0 PWL(0 0 'input_delay3+0*trf_ip_reset+0*input_pw' 0 'input_delay3+1*trf_ip_reset+0*input_pw' 0 'input_delay3+1*trf_ip_reset+1*input_pw' 0 'input_delay3+2*trf_ip_reset+1*input_pw' 0 'input_delay3+2*trf_ip_reset+2*input_pw' 0 'input_delay3+3*trf_ip_reset+2*input_pw' 1.8 'input_delay3+3*trf_ip_reset+3*input_pw' 1.8  'input_delay3+4*trf_ip_reset+3*input_pw' 0 'input_delay3+4*trf_ip_reset+4*input_pw' 0 'input_delay3+5*trf_ip_reset+4*input_pw' 1.8 sim_end 1.8)
vA1 a1 0 PWL(0 0 'input_delay4+0*trf_ip_reset+0*input_pw' 0 'input_delay4+1*trf_ip_reset+0*input_pw' 1.8 'input_delay4+1*trf_ip_reset+1*input_pw' 1.8 'input_delay4+2*trf_ip_reset+1*input_pw' 1.8 'input_delay4+2*trf_ip_reset+2*input_pw' 1.8 'input_delay4+3*trf_ip_reset+2*input_pw' 1.8 'input_delay4+3*trf_ip_reset+3*input_pw' 1.8  'input_delay4+4*trf_ip_reset+3*input_pw' 1.8 'input_delay4+4*trf_ip_reset+4*input_pw' 1.8 'input_delay4+5*trf_ip_reset+4*input_pw' 0 sim_end 0)
vB3 b3 0 PWL(0 0 'input_delay2+0*trf_ip_reset+0*input_pw' 0 'input_delay2+1*trf_ip_reset+0*input_pw' 1.8 'input_delay2+1*trf_ip_reset+1*input_pw' 1.8 'input_delay2+2*trf_ip_reset+1*input_pw' 1.8 'input_delay2+2*trf_ip_reset+2*input_pw' 1.8 'input_delay2+3*trf_ip_reset+2*input_pw' 1.8 'input_delay2+3*trf_ip_reset+3*input_pw' 1.8  'input_delay2+4*trf_ip_reset+3*input_pw' 0 'input_delay2+4*trf_ip_reset+4*input_pw' 0 'input_delay2+5*trf_ip_reset+4*input_pw' 1.8 sim_end 1.8)
vB1 b1 0 PWL(0 0 'input_delay+0*trf_ip_reset+0*input_pw' 0 'input_delay+1*trf_ip_reset+0*input_pw' 0 'input_delay+1*trf_ip_reset+1*input_pw' 0 'input_delay+2*trf_ip_reset+1*input_pw' 0 'input_delay+2*trf_ip_reset+2*input_pw' 0 'input_delay+2*trf_ip_reset+2*input_pw+offset_ip' 0 'input_delay+3*trf_ip_reset+2*input_pw+offset_ip' 1.8 'input_delay+3*trf_ip_reset+3*input_pw+offset_ip' 1.8  'input_delay+4*trf_ip_reset+3*input_pw+offset_ip' 1.8 'input_delay+4*trf_ip_reset+4*input_pw+offset_ip' 1.8 'input_delay+5*trf_ip_reset+4*input_pw+offset_ip' 1.8 sim_end 1.8)
vB0 b0 0 PWL(0 0 'input_delay2+0*trf_ip_reset+0*input_pw' 0 'input_delay2+1*trf_ip_reset+0*input_pw' 0 'input_delay2+1*trf_ip_reset+1*input_pw' 0 'input_delay2+2*trf_ip_reset+1*input_pw' 1.8 'input_delay2+2*trf_ip_reset+2*input_pw' 1.8 'input_delay2+3*trf_ip_reset+2*input_pw' 1.8 'input_delay2+3*trf_ip_reset+3*input_pw' 1.8  'input_delay2+4*trf_ip_reset+3*input_pw' 0 'input_delay2+4*trf_ip_reset+4*input_pw' 0 'input_delay2+5*trf_ip_reset+4*input_pw' 1.8 sim_end 1.8)
vB2 b2 0 PWL(0 0 'input_delay4+0*trf_ip_reset+0*input_pw' 0 'input_delay4+1*trf_ip_reset+0*input_pw' 0 'input_delay4+1*trf_ip_reset+1*input_pw' 0 'input_delay4+2*trf_ip_reset+1*input_pw' 0 'input_delay4+2*trf_ip_reset+2*input_pw' 0 'input_delay4+3*trf_ip_reset+2*input_pw' 1.8 'input_delay4+3*trf_ip_reset+3*input_pw' 1.8  'input_delay4+4*trf_ip_reset+3*input_pw' 1.8 'input_delay4+4*trf_ip_reset+4*input_pw' 1.8 'input_delay4+5*trf_ip_reset+4*input_pw' 1.8 sim_end 1.8)

*Sources on board - ONly nom_vdd value can be modified for power reduction using the parameters above.
vVDDIO VDDIO 0 1.8
vVDD VDD 0 nom_vdd
vVSS VSS 0 0

*Bondwire inductance - Not to be modified.
LVSS1 vss1 VSS 2.5n
LVSS2 vss2 VSS 2.5n
LVSS3 vss3 VSS 2.5n
LVSS4 vss4 VSS 2.5n
LVSSIO1 vssio1 VSS 2.5n
LVSSIO2 vssio2 VSS 2.5n
LVSSIO3 vssio3 VSS 2.5n
LVDDIO1 vddio1 VDDIO 5n
LVDDIO2 vddio2 VDDIO 5n
LVDDIO3 vddio3 VDDIO 5n
LVDD1 vdd1 VDD 5n
LVDD2 vdd2 VDD 5n
LVDD3 vdd3 VDD 5n

LA0 a0 a0_oc 4n
LA1 a1 a1_oc 4n
LA2 a2 a2_oc 4n
LA3 a3 a3_oc 4n
LB0 b0 b0_oc 4n
LB1 b1 b1_oc 4n
LB2 b2 b2_oc 4n
LB3 b3 b3_oc 4n

LP0 p0 p0_oc 4n
LP1 p1 p1_oc 4n
LP2 p2 p2_oc 4n
LP3 p3 p3_oc 4n
LP4 p4 p4_oc 4n
LP5 p5 p5_oc 4n
LP6 p6 p6_oc 4n
LP7 p7 p7_oc 4n

LRST reset rst_oc 4n
LCLK clk clk_oc 2n

*ESD capacitance - Not to be modified.
CVDD1 vdd1 vss1 0.3p
CVDD2 vdd2 vss2 0.3p
CVDD3 vdd3 vss3 0.3p
CVDDIO1 vdd1 vss1 0.4p
CVDDIO2 vdd2 vss2 0.4p
CVDDIO3 vdd3 vss3 0.4p

CA0_OC a0_oc1 vss4 0.25p
CA1_OC a1_oc1 vssio1 0.25p
CA2_OC a2_oc1 vssio2 0.25p
CA3_OC a3_oc1 vssio3 0.25p
CB0_OC b0_oc1 vss1 0.25p
CB1_OC b1_oc1 vss2 0.25p
CB2_OC b2_oc1 vss3 0.25p
CB3_OC b3_oc1 vss4 0.25p

CP0_OC p0_oc1 vss4 0.25p
CP1_OC p1_oc1 vssio1 0.25p
CP2_OC p2_oc1 vssio2 0.25p
CP3_OC p3_oc1 vssio3 0.25p
CP4_OC p4_oc1 vss1 0.25p
CP5_OC p5_oc1 vss2 0.25p
CP6_OC p6_oc1 vss3 0.25p
CP7_OC p7_oc1 vss4 0.25p


CCLK_OC clk_oc1 vss1 0.3p
CRST_OC rst_oc1 vss1 0.25p

*Load Capacitance - Not to be modified.
CA0 a0 VSS 20p
CA1 a1 VSS 20p
CA2 a2 VSS 20p
CA3 a3 VSS 20p
CB0 b0 VSS 20p
CB1 b1 VSS 20p
CB2 b2 VSS 20p
CB3 b3 VSS 20p

CP0 p0 VSS 20p
CP1 p1 VSS 20p
CP2 p2 VSS 20p
CP3 p3 VSS 20p
CP4 p4 VSS 20p
CP5 p5 VSS 20p
CP6 p6 VSS 20p
CP7 p7 VSS 20p


CCLK clk VSS 2p
CRST reset VSS 20p

.tran 0 sim_end

*Power measurement functions - NOt to be modified.
.meas tran avg_pwr_vdd avg p(vVDD) from=reset_delay+reset_pw+2*trf_ip_reset to=sim_end-2n
.meas tran avg_pwr_vddio avg p(vVDDIO) from=reset_delay+reset_pw+2*trf_ip_reset to=sim_end-2n
* Corrected power after subtracting noisy current source power
.meas tran corrected_pwr_vdd  param='avg_pwr_vdd + 0.0217681251338'

.probe tran i(ILOAD)
.print tran vdd_net='v(vdd1) - v(vss1)'
.print tran vddio_net='v(vddio1) - v(vssio1)'
.option post
.end
